`include "define.v"                                       
 module R16_WD_buf(RDC0_D_out,                               
 			       RDC1_D_out,                              
 				   RDC2_D_out,                              
 				   RDC3_D_out,                              
 				   RDC4_D_out,                              
 				   RDC5_D_out,                              
 				   RDC6_D_out,                              
 				   RDC7_D_out,                              
 				   RDC8_D_out,                              
 				   RDC9_D_out,                              
 				   RDC10_D_out,                             
 				   RDC11_D_out,                             
 				   RDC12_D_out,                             
 				   RDC13_D_out,                             
 				   RDC14_D_out,                             
 				   RDC15_D_out,                             
 		           RDC0_in,                                 
 				   RDC1_in,                                 
 				   RDC2_in,                                 
 				   RDC3_in,                                 
 				   RDC4_in,                                 
 				   RDC5_in,                                 
 				   RDC6_in,                                 
 				   RDC7_in,                                 
 				   RDC8_in,                                 
 				   RDC9_in,                                 
 				   RDC10_in,                                
 				   RDC11_in,                                
 				   RDC12_in,                                
 				   RDC13_in,                                
 				   RDC14_in,                                
 				   RDC15_in,                                
                   rst_n,                                    
                   clk                                       
                   ) ;                                       
 parameter P_WIDTH     = 64 ;                                
                                                             
 parameter P_ZERO    = 64'h0 ;                               
                                                             
                                                             
 output [P_WIDTH-1:0] RDC0_D_out ;                           
 output [P_WIDTH-1:0] RDC1_D_out ;                           
 output [P_WIDTH-1:0] RDC2_D_out ;                           
 output [P_WIDTH-1:0] RDC3_D_out ;                           
 output [P_WIDTH-1:0] RDC4_D_out ;                           
 output [P_WIDTH-1:0] RDC5_D_out ;                           
 output [P_WIDTH-1:0] RDC6_D_out ;                           
 output [P_WIDTH-1:0] RDC7_D_out ;                           
 output [P_WIDTH-1:0] RDC8_D_out ;                           
 output [P_WIDTH-1:0] RDC9_D_out ;                           
 output [P_WIDTH-1:0] RDC10_D_out ;                          
 output [P_WIDTH-1:0] RDC11_D_out ;                          
 output [P_WIDTH-1:0] RDC12_D_out ;                          
 output [P_WIDTH-1:0] RDC13_D_out ;                          
 output [P_WIDTH-1:0] RDC14_D_out ;                          
 output [P_WIDTH-1:0] RDC15_D_out ;                          
                                                             
 input [P_WIDTH-1:0] RDC0_in ;                               
 input [P_WIDTH-1:0] RDC1_in ;                               
 input [P_WIDTH-1:0] RDC2_in ;                               
 input [P_WIDTH-1:0] RDC3_in ;                               
 input [P_WIDTH-1:0] RDC4_in ;                               
 input [P_WIDTH-1:0] RDC5_in ;                               
 input [P_WIDTH-1:0] RDC6_in ;                               
 input [P_WIDTH-1:0] RDC7_in ;                               
 input [P_WIDTH-1:0] RDC8_in ;                               
 input [P_WIDTH-1:0] RDC9_in ;                               
 input [P_WIDTH-1:0] RDC10_in ;                              
 input [P_WIDTH-1:0] RDC11_in ;                              
 input [P_WIDTH-1:0] RDC12_in ;                              
 input [P_WIDTH-1:0] RDC13_in ;                              
 input [P_WIDTH-1:0] RDC14_in ;                              
 input [P_WIDTH-1:0] RDC15_in ;                              
 input               rst_n ;                                 
 input               clk ;                                   
                                                             
                                                             
 reg  [P_WIDTH-1:0] RDC0_D_out ;                             
 reg  [P_WIDTH-1:0] RDC1_D_out ;                             
 reg  [P_WIDTH-1:0] RDC2_D_out ;                             
 reg  [P_WIDTH-1:0] RDC3_D_out ;                             
 reg  [P_WIDTH-1:0] RDC4_D_out ;                             
 reg  [P_WIDTH-1:0] RDC5_D_out ;                             
 reg  [P_WIDTH-1:0] RDC6_D_out ;                             
 reg  [P_WIDTH-1:0] RDC7_D_out ;                             
 reg  [P_WIDTH-1:0] RDC8_D_out ;                             
 reg  [P_WIDTH-1:0] RDC9_D_out ;                             
 reg  [P_WIDTH-1:0] RDC10_D_out ;                            
 reg  [P_WIDTH-1:0] RDC11_D_out ;                            
 reg  [P_WIDTH-1:0] RDC12_D_out ;                            
 reg  [P_WIDTH-1:0] RDC13_D_out ;                            
 reg  [P_WIDTH-1:0] RDC14_D_out ;                            
 reg  [P_WIDTH-1:0] RDC15_D_out ;                            
                                                             
 reg  [P_WIDTH-1:0] RDC0_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC0_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC0_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC0_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC1_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC1_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC1_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC1_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC2_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC2_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC2_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC2_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC3_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC3_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC3_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC3_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC4_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC4_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC4_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC4_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC5_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC5_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC5_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC5_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC6_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC6_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC6_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC6_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC7_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC7_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC7_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC7_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC8_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC8_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC8_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC8_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC9_D0_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D1_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D2_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D3_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D4_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D5_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D6_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D7_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D8_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D9_reg ;                            
 reg  [P_WIDTH-1:0] RDC9_D10_reg ;                           
 reg  [P_WIDTH-1:0] RDC9_D11_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D12_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D13_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D14_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D15_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D16_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D17_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D18_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D19_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D20_reg  ;                          
 reg  [P_WIDTH-1:0] RDC9_D21_reg  ;                          
                                                             
 reg  [P_WIDTH-1:0] RDC10_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC10_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC10_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC10_D21_reg  ;                         
                                                             
 reg  [P_WIDTH-1:0] RDC11_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC11_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC11_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC11_D21_reg  ;                         
                                                             
 reg  [P_WIDTH-1:0] RDC12_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC12_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC12_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC12_D21_reg  ;                         
                                                             
 reg  [P_WIDTH-1:0] RDC13_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC13_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC13_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC13_D21_reg  ;                         
                                                             
 reg  [P_WIDTH-1:0] RDC14_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC14_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC14_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC14_D21_reg  ;                         
                                                             
 reg  [P_WIDTH-1:0] RDC15_D0_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D1_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D2_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D3_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D4_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D5_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D6_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D7_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D8_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D9_reg ;                           
 reg  [P_WIDTH-1:0] RDC15_D10_reg ;                          
 reg  [P_WIDTH-1:0] RDC15_D11_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D12_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D13_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D14_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D15_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D16_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D17_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D18_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D19_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D20_reg  ;                         
 reg  [P_WIDTH-1:0] RDC15_D21_reg  ;                         
                                                             
 	//RDC output delay 23 cycles                            
 	always @(posedge clk or negedge rst_n) begin            
 		if(~rst_n) begin                                    
 			RDC0_D0_reg  <= P_ZERO ;                        
 			RDC0_D1_reg  <= P_ZERO;                         
 			RDC0_D2_reg  <= P_ZERO;                         
 			RDC0_D3_reg  <= P_ZERO;                         
 			RDC0_D4_reg  <= P_ZERO;                         
 			RDC0_D5_reg  <= P_ZERO;                         
 			RDC0_D6_reg  <= P_ZERO;                         
 			RDC0_D7_reg  <= P_ZERO;                         
 			RDC0_D8_reg  <= P_ZERO;                         
 			RDC0_D9_reg  <= P_ZERO;                         
 			RDC0_D10_reg <= P_ZERO;                         
 			RDC0_D11_reg <= P_ZERO ;                        
 			RDC0_D12_reg <= P_ZERO ;                        
 			RDC0_D13_reg <= P_ZERO ;                        
 			RDC0_D14_reg <= P_ZERO ;                        
 			RDC0_D15_reg <= P_ZERO ;                        
 			RDC0_D16_reg <= P_ZERO ;                        
 			RDC0_D17_reg <= P_ZERO ;                        
 			RDC0_D18_reg <= P_ZERO ;                        
 			RDC0_D19_reg <= P_ZERO ;                        
 			RDC0_D20_reg <= P_ZERO ;                        
 			RDC0_D21_reg <= P_ZERO ;                        
 			RDC0_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC1_D0_reg  <= P_ZERO ;                        
 			RDC1_D1_reg  <= P_ZERO;                         
 			RDC1_D2_reg  <= P_ZERO;                         
 			RDC1_D3_reg  <= P_ZERO;                         
 			RDC1_D4_reg  <= P_ZERO;                         
 			RDC1_D5_reg  <= P_ZERO;                         
 			RDC1_D6_reg  <= P_ZERO;                         
 			RDC1_D7_reg  <= P_ZERO;                         
 			RDC1_D8_reg  <= P_ZERO;                         
 			RDC1_D9_reg  <= P_ZERO;                         
 			RDC1_D10_reg <= P_ZERO;                         
 			RDC1_D11_reg <= P_ZERO ;                        
 			RDC1_D12_reg <= P_ZERO ;                        
 			RDC1_D13_reg <= P_ZERO ;                        
 			RDC1_D14_reg <= P_ZERO ;                        
 			RDC1_D15_reg <= P_ZERO ;                        
 			RDC1_D16_reg <= P_ZERO ;                        
 			RDC1_D17_reg <= P_ZERO ;                        
 			RDC1_D18_reg <= P_ZERO ;                        
 			RDC1_D19_reg <= P_ZERO ;                        
 			RDC1_D20_reg <= P_ZERO ;                        
 			RDC1_D21_reg <= P_ZERO ;                        
 			RDC1_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC2_D0_reg  <= P_ZERO ;                        
 			RDC2_D1_reg  <= P_ZERO;                         
 			RDC2_D2_reg  <= P_ZERO;                         
 			RDC2_D3_reg  <= P_ZERO;                         
 			RDC2_D4_reg  <= P_ZERO;                         
 			RDC2_D5_reg  <= P_ZERO;                         
 			RDC2_D6_reg  <= P_ZERO;                         
 			RDC2_D7_reg  <= P_ZERO;                         
 			RDC2_D8_reg  <= P_ZERO;                         
 			RDC2_D9_reg  <= P_ZERO;                         
 			RDC2_D10_reg <= P_ZERO;                         
 			RDC2_D11_reg <= P_ZERO ;                        
 			RDC2_D12_reg <= P_ZERO ;                        
 			RDC2_D13_reg <= P_ZERO ;                        
 			RDC2_D14_reg <= P_ZERO ;                        
 			RDC2_D15_reg <= P_ZERO ;                        
 			RDC2_D16_reg <= P_ZERO ;                        
 			RDC2_D17_reg <= P_ZERO ;                        
 			RDC2_D18_reg <= P_ZERO ;                        
 			RDC2_D19_reg <= P_ZERO ;                        
 			RDC2_D20_reg <= P_ZERO ;                        
 			RDC2_D21_reg <= P_ZERO ;                        
 			RDC2_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC3_D0_reg  <= P_ZERO ;                        
 			RDC3_D1_reg  <= P_ZERO;                         
 			RDC3_D2_reg  <= P_ZERO;                         
 			RDC3_D3_reg  <= P_ZERO;                         
 			RDC3_D4_reg  <= P_ZERO;                         
 			RDC3_D5_reg  <= P_ZERO;                         
 			RDC3_D6_reg  <= P_ZERO;                         
 			RDC3_D7_reg  <= P_ZERO;                         
 			RDC3_D8_reg  <= P_ZERO;                         
 			RDC3_D9_reg  <= P_ZERO;                         
 			RDC3_D10_reg <= P_ZERO;                         
 			RDC3_D11_reg <= P_ZERO ;                        
 			RDC3_D12_reg <= P_ZERO ;                        
 			RDC3_D13_reg <= P_ZERO ;                        
 			RDC3_D14_reg <= P_ZERO ;                        
 			RDC3_D15_reg <= P_ZERO ;                        
 			RDC3_D16_reg <= P_ZERO ;                        
 			RDC3_D17_reg <= P_ZERO ;                        
 			RDC3_D18_reg <= P_ZERO ;                        
 			RDC3_D19_reg <= P_ZERO ;                        
 			RDC3_D20_reg <= P_ZERO ;                        
 			RDC3_D21_reg <= P_ZERO ;                        
 			RDC3_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC4_D0_reg  <= P_ZERO ;                        
 			RDC4_D1_reg  <= P_ZERO;                         
 			RDC4_D2_reg  <= P_ZERO;                         
 			RDC4_D3_reg  <= P_ZERO;                         
 			RDC4_D4_reg  <= P_ZERO;                         
 			RDC4_D5_reg  <= P_ZERO;                         
 			RDC4_D6_reg  <= P_ZERO;                         
 			RDC4_D7_reg  <= P_ZERO;                         
 			RDC4_D8_reg  <= P_ZERO;                         
 			RDC4_D9_reg  <= P_ZERO;                         
 			RDC4_D10_reg <= P_ZERO;                         
 			RDC4_D11_reg <= P_ZERO ;                        
 			RDC4_D12_reg <= P_ZERO ;                        
 			RDC4_D13_reg <= P_ZERO ;                        
 			RDC4_D14_reg <= P_ZERO ;                        
 			RDC4_D15_reg <= P_ZERO ;                        
 			RDC4_D16_reg <= P_ZERO ;                        
 			RDC4_D17_reg <= P_ZERO ;                        
 			RDC4_D18_reg <= P_ZERO ;                        
 			RDC4_D19_reg <= P_ZERO ;                        
 			RDC4_D20_reg <= P_ZERO ;                        
 			RDC4_D21_reg <= P_ZERO ;                        
 			RDC4_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC5_D0_reg  <= P_ZERO ;                        
 			RDC5_D1_reg  <= P_ZERO;                         
 			RDC5_D2_reg  <= P_ZERO;                         
 			RDC5_D3_reg  <= P_ZERO;                         
 			RDC5_D4_reg  <= P_ZERO;                         
 			RDC5_D5_reg  <= P_ZERO;                         
 			RDC5_D6_reg  <= P_ZERO;                         
 			RDC5_D7_reg  <= P_ZERO;                         
 			RDC5_D8_reg  <= P_ZERO;                         
 			RDC5_D9_reg  <= P_ZERO;                         
 			RDC5_D10_reg <= P_ZERO;                         
 			RDC5_D11_reg <= P_ZERO ;                        
 			RDC5_D12_reg <= P_ZERO ;                        
 			RDC5_D13_reg <= P_ZERO ;                        
 			RDC5_D14_reg <= P_ZERO ;                        
 			RDC5_D15_reg <= P_ZERO ;                        
 			RDC5_D16_reg <= P_ZERO ;                        
 			RDC5_D17_reg <= P_ZERO ;                        
 			RDC5_D18_reg <= P_ZERO ;                        
 			RDC5_D19_reg <= P_ZERO ;                        
 			RDC5_D20_reg <= P_ZERO ;                        
 			RDC5_D21_reg <= P_ZERO ;                        
 			RDC5_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC6_D0_reg  <= P_ZERO ;                        
 			RDC6_D1_reg  <= P_ZERO;                         
 			RDC6_D2_reg  <= P_ZERO;                         
 			RDC6_D3_reg  <= P_ZERO;                         
 			RDC6_D4_reg  <= P_ZERO;                         
 			RDC6_D5_reg  <= P_ZERO;                         
 			RDC6_D6_reg  <= P_ZERO;                         
 			RDC6_D7_reg  <= P_ZERO;                         
 			RDC6_D8_reg  <= P_ZERO;                         
 			RDC6_D9_reg  <= P_ZERO;                         
 			RDC6_D10_reg <= P_ZERO;                         
 			RDC6_D11_reg <= P_ZERO ;                        
 			RDC6_D12_reg <= P_ZERO ;                        
 			RDC6_D13_reg <= P_ZERO ;                        
 			RDC6_D14_reg <= P_ZERO ;                        
 			RDC6_D15_reg <= P_ZERO ;                        
 			RDC6_D16_reg <= P_ZERO ;                        
 			RDC6_D17_reg <= P_ZERO ;                        
 			RDC6_D18_reg <= P_ZERO ;                        
 			RDC6_D19_reg <= P_ZERO ;                        
 			RDC6_D20_reg <= P_ZERO ;                        
 			RDC6_D21_reg <= P_ZERO ;                        
 			RDC6_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC7_D0_reg  <= P_ZERO ;                        
 			RDC7_D1_reg  <= P_ZERO;                         
 			RDC7_D2_reg  <= P_ZERO;                         
 			RDC7_D3_reg  <= P_ZERO;                         
 			RDC7_D4_reg  <= P_ZERO;                         
 			RDC7_D5_reg  <= P_ZERO;                         
 			RDC7_D6_reg  <= P_ZERO;                         
 			RDC7_D7_reg  <= P_ZERO;                         
 			RDC7_D8_reg  <= P_ZERO;                         
 			RDC7_D9_reg  <= P_ZERO;                         
 			RDC7_D10_reg <= P_ZERO;                         
 			RDC7_D11_reg <= P_ZERO ;                        
 			RDC7_D12_reg <= P_ZERO ;                        
 			RDC7_D13_reg <= P_ZERO ;                        
 			RDC7_D14_reg <= P_ZERO ;                        
 			RDC7_D15_reg <= P_ZERO ;                        
 			RDC7_D16_reg <= P_ZERO ;                        
 			RDC7_D17_reg <= P_ZERO ;                        
 			RDC7_D18_reg <= P_ZERO ;                        
 			RDC7_D19_reg <= P_ZERO ;                        
 			RDC7_D20_reg <= P_ZERO ;                        
 			RDC7_D21_reg <= P_ZERO ;                        
 			RDC7_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC8_D0_reg  <= P_ZERO ;                        
 			RDC8_D1_reg  <= P_ZERO;                         
 			RDC8_D2_reg  <= P_ZERO;                         
 			RDC8_D3_reg  <= P_ZERO;                         
 			RDC8_D4_reg  <= P_ZERO;                         
 			RDC8_D5_reg  <= P_ZERO;                         
 			RDC8_D6_reg  <= P_ZERO;                         
 			RDC8_D7_reg  <= P_ZERO;                         
 			RDC8_D8_reg  <= P_ZERO;                         
 			RDC8_D9_reg  <= P_ZERO;                         
 			RDC8_D10_reg <= P_ZERO;                         
 			RDC8_D11_reg <= P_ZERO ;                        
 			RDC8_D12_reg <= P_ZERO ;                        
 			RDC8_D13_reg <= P_ZERO ;                        
 			RDC8_D14_reg <= P_ZERO ;                        
 			RDC8_D15_reg <= P_ZERO ;                        
 			RDC8_D16_reg <= P_ZERO ;                        
 			RDC8_D17_reg <= P_ZERO ;                        
 			RDC8_D18_reg <= P_ZERO ;                        
 			RDC8_D19_reg <= P_ZERO ;                        
 			RDC8_D20_reg <= P_ZERO ;                        
 			RDC8_D21_reg <= P_ZERO ;                        
 			RDC8_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC9_D0_reg  <= P_ZERO ;                        
 			RDC9_D1_reg  <= P_ZERO;                         
 			RDC9_D2_reg  <= P_ZERO;                         
 			RDC9_D3_reg  <= P_ZERO;                         
 			RDC9_D4_reg  <= P_ZERO;                         
 			RDC9_D5_reg  <= P_ZERO;                         
 			RDC9_D6_reg  <= P_ZERO;                         
 			RDC9_D7_reg  <= P_ZERO;                         
 			RDC9_D8_reg  <= P_ZERO;                         
 			RDC9_D9_reg  <= P_ZERO;                         
 			RDC9_D10_reg <= P_ZERO;                         
 			RDC9_D11_reg <= P_ZERO ;                        
 			RDC9_D12_reg <= P_ZERO ;                        
 			RDC9_D13_reg <= P_ZERO ;                        
 			RDC9_D14_reg <= P_ZERO ;                        
 			RDC9_D15_reg <= P_ZERO ;                        
 			RDC9_D16_reg <= P_ZERO ;                        
 			RDC9_D17_reg <= P_ZERO ;                        
 			RDC9_D18_reg <= P_ZERO ;                        
 			RDC9_D19_reg <= P_ZERO ;                        
 			RDC9_D20_reg <= P_ZERO ;                        
 			RDC9_D21_reg <= P_ZERO ;                        
 			RDC9_D_out   <= P_ZERO ;                        
 			//                                              
 			RDC10_D0_reg  <= P_ZERO ;                       
 			RDC10_D1_reg  <= P_ZERO;                        
 			RDC10_D2_reg  <= P_ZERO;                        
 			RDC10_D3_reg  <= P_ZERO;                        
 			RDC10_D4_reg  <= P_ZERO;                        
 			RDC10_D5_reg  <= P_ZERO;                        
 			RDC10_D6_reg  <= P_ZERO;                        
 			RDC10_D7_reg  <= P_ZERO;                        
 			RDC10_D8_reg  <= P_ZERO;                        
 			RDC10_D9_reg  <= P_ZERO;                        
 			RDC10_D10_reg <= P_ZERO;                        
 			RDC10_D11_reg <= P_ZERO ;                       
 			RDC10_D12_reg <= P_ZERO ;                       
 			RDC10_D13_reg <= P_ZERO ;                       
 			RDC10_D14_reg <= P_ZERO ;                       
 			RDC10_D15_reg <= P_ZERO ;                       
 			RDC10_D16_reg <= P_ZERO ;                       
 			RDC10_D17_reg <= P_ZERO ;                       
 			RDC10_D18_reg <= P_ZERO ;                       
 			RDC10_D19_reg <= P_ZERO ;                       
 			RDC10_D20_reg <= P_ZERO ;                       
 			RDC10_D21_reg <= P_ZERO ;                       
 			RDC10_D_out   <= P_ZERO ;                       
 			//                                              
 			RDC11_D0_reg  <= P_ZERO ;                       
 			RDC11_D1_reg  <= P_ZERO;                        
 			RDC11_D2_reg  <= P_ZERO;                        
 			RDC11_D3_reg  <= P_ZERO;                        
 			RDC11_D4_reg  <= P_ZERO;                        
 			RDC11_D5_reg  <= P_ZERO;                        
 			RDC11_D6_reg  <= P_ZERO;                        
 			RDC11_D7_reg  <= P_ZERO;                        
 			RDC11_D8_reg  <= P_ZERO;                        
 			RDC11_D9_reg  <= P_ZERO;                        
 			RDC11_D10_reg <= P_ZERO;                        
 			RDC11_D11_reg <= P_ZERO ;                       
 			RDC11_D12_reg <= P_ZERO ;                       
 			RDC11_D13_reg <= P_ZERO ;                       
 			RDC11_D14_reg <= P_ZERO ;                       
 			RDC11_D15_reg <= P_ZERO ;                       
 			RDC11_D16_reg <= P_ZERO ;                       
 			RDC11_D17_reg <= P_ZERO ;                       
 			RDC11_D18_reg <= P_ZERO ;                       
 			RDC11_D19_reg <= P_ZERO ;                       
 			RDC11_D20_reg <= P_ZERO ;                       
 			RDC11_D21_reg <= P_ZERO ;                       
 			RDC11_D_out   <= P_ZERO ;                       
 			//                                              
 			RDC12_D0_reg  <= P_ZERO ;                       
 			RDC12_D1_reg  <= P_ZERO;                        
 			RDC12_D2_reg  <= P_ZERO;                        
 			RDC12_D3_reg  <= P_ZERO;                        
 			RDC12_D4_reg  <= P_ZERO;                        
 			RDC12_D5_reg  <= P_ZERO;                        
 			RDC12_D6_reg  <= P_ZERO;                        
 			RDC12_D7_reg  <= P_ZERO;                        
 			RDC12_D8_reg  <= P_ZERO;                        
 			RDC12_D9_reg  <= P_ZERO;                        
 			RDC12_D10_reg <= P_ZERO;                        
 			RDC12_D11_reg <= P_ZERO ;                       
 			RDC12_D12_reg <= P_ZERO ;                       
 			RDC12_D13_reg <= P_ZERO ;                       
 			RDC12_D14_reg <= P_ZERO ;                       
 			RDC12_D15_reg <= P_ZERO ;                       
 			RDC12_D16_reg <= P_ZERO ;                       
 			RDC12_D17_reg <= P_ZERO ;                       
 			RDC12_D18_reg <= P_ZERO ;                       
 			RDC12_D19_reg <= P_ZERO ;                       
 			RDC12_D20_reg <= P_ZERO ;                       
 			RDC12_D21_reg <= P_ZERO ;                       
 			RDC12_D_out   <= P_ZERO ;                       
 			//                                              
 			RDC13_D0_reg  <= P_ZERO ;                       
 			RDC13_D1_reg  <= P_ZERO;                        
 			RDC13_D2_reg  <= P_ZERO;                        
 			RDC13_D3_reg  <= P_ZERO;                        
 			RDC13_D4_reg  <= P_ZERO;                        
 			RDC13_D5_reg  <= P_ZERO;                        
 			RDC13_D6_reg  <= P_ZERO;                        
 			RDC13_D7_reg  <= P_ZERO;                        
 			RDC13_D8_reg  <= P_ZERO;                        
 			RDC13_D9_reg  <= P_ZERO;                        
 			RDC13_D10_reg <= P_ZERO;                        
 			RDC13_D11_reg <= P_ZERO ;                       
 			RDC13_D12_reg <= P_ZERO ;                       
 			RDC13_D13_reg <= P_ZERO ;                       
 			RDC13_D14_reg <= P_ZERO ;                       
 			RDC13_D15_reg <= P_ZERO ;                       
 			RDC13_D16_reg <= P_ZERO ;                       
 			RDC13_D17_reg <= P_ZERO ;                       
 			RDC13_D18_reg <= P_ZERO ;                       
 			RDC13_D19_reg <= P_ZERO ;                       
 			RDC13_D20_reg <= P_ZERO ;                       
 			RDC13_D21_reg <= P_ZERO ;                       
 			RDC13_D_out   <= P_ZERO ;                       
 			//                                              
 			RDC14_D0_reg  <= P_ZERO ;                       
 			RDC14_D1_reg  <= P_ZERO;                        
 			RDC14_D2_reg  <= P_ZERO;                        
 			RDC14_D3_reg  <= P_ZERO;                        
 			RDC14_D4_reg  <= P_ZERO;                        
 			RDC14_D5_reg  <= P_ZERO;                        
 			RDC14_D6_reg  <= P_ZERO;                        
 			RDC14_D7_reg  <= P_ZERO;                        
 			RDC14_D8_reg  <= P_ZERO;                        
 			RDC14_D9_reg  <= P_ZERO;                        
 			RDC14_D10_reg <= P_ZERO;                        
 			RDC14_D11_reg <= P_ZERO ;                       
 			RDC14_D12_reg <= P_ZERO ;                       
 			RDC14_D13_reg <= P_ZERO ;                       
 			RDC14_D14_reg <= P_ZERO ;                       
 			RDC14_D15_reg <= P_ZERO ;                       
 			RDC14_D16_reg <= P_ZERO ;                       
 			RDC14_D17_reg <= P_ZERO ;                       
 			RDC14_D18_reg <= P_ZERO ;                       
 			RDC14_D19_reg <= P_ZERO ;                       
 			RDC14_D20_reg <= P_ZERO ;                       
 			RDC14_D21_reg <= P_ZERO ;                       
 			RDC14_D_out   <= P_ZERO ;                       
 			//                                              
 			RDC15_D0_reg  <= P_ZERO ;                       
 			RDC15_D1_reg  <= P_ZERO;                        
 			RDC15_D2_reg  <= P_ZERO;                        
 			RDC15_D3_reg  <= P_ZERO;                        
 			RDC15_D4_reg  <= P_ZERO;                        
 			RDC15_D5_reg  <= P_ZERO;                        
 			RDC15_D6_reg  <= P_ZERO;                        
 			RDC15_D7_reg  <= P_ZERO;                        
 			RDC15_D8_reg  <= P_ZERO;                        
 			RDC15_D9_reg  <= P_ZERO;                        
 			RDC15_D10_reg <= P_ZERO;                        
 			RDC15_D11_reg <= P_ZERO ;                       
 			RDC15_D12_reg <= P_ZERO ;                       
 			RDC15_D13_reg <= P_ZERO ;                       
 			RDC15_D14_reg <= P_ZERO ;                       
 			RDC15_D15_reg <= P_ZERO ;                       
 			RDC15_D16_reg <= P_ZERO ;                       
 			RDC15_D17_reg <= P_ZERO ;                       
 			RDC15_D18_reg <= P_ZERO ;                       
 			RDC15_D19_reg <= P_ZERO ;                       
 			RDC15_D20_reg <= P_ZERO ;                       
 			RDC15_D21_reg <= P_ZERO ;                       
 			RDC15_D_out   <= P_ZERO ;                       
 		end                                                 
 		else begin                                          
 			RDC0_D0_reg  <= RDC0_in ;                       
 			RDC0_D1_reg  <= RDC0_D0_reg ;                   
 			RDC0_D2_reg  <= RDC0_D1_reg ;                   
 			RDC0_D3_reg  <= RDC0_D2_reg ;                   
 			RDC0_D4_reg  <= RDC0_D3_reg ;                   
 			RDC0_D5_reg  <= RDC0_D4_reg ;                   
 			RDC0_D6_reg  <= RDC0_D5_reg ;                   
 			RDC0_D7_reg  <= RDC0_D6_reg ;                   
 			RDC0_D8_reg  <= RDC0_D7_reg ;                   
 			RDC0_D9_reg  <= RDC0_D8_reg ;                   
 			RDC0_D10_reg <= RDC0_D9_reg ;                   
 			RDC0_D11_reg <= RDC0_D10_reg ;                  
 			RDC0_D12_reg <= RDC0_D11_reg ;                  
 			RDC0_D13_reg <= RDC0_D12_reg ;                  
 			RDC0_D14_reg <= RDC0_D13_reg ;                  
 			RDC0_D15_reg <= RDC0_D14_reg ;                  
 			RDC0_D16_reg <= RDC0_D15_reg ;                  
 			RDC0_D17_reg <= RDC0_D16_reg ;                  
 			RDC0_D18_reg <= RDC0_D17_reg ;                  
 			RDC0_D19_reg <= RDC0_D18_reg ;                  
 			RDC0_D20_reg <= RDC0_D19_reg ;                  
 			RDC0_D21_reg <= RDC0_D20_reg ;                  
 			RDC0_D_out   <= RDC0_D21_reg ;                  
 			//                                              
 			RDC1_D0_reg  <= RDC1_in ;                       
 			RDC1_D1_reg  <= RDC1_D0_reg ;                   
 			RDC1_D2_reg  <= RDC1_D1_reg ;                   
 			RDC1_D3_reg  <= RDC1_D2_reg ;                   
 			RDC1_D4_reg  <= RDC1_D3_reg ;                   
 			RDC1_D5_reg  <= RDC1_D4_reg ;                   
 			RDC1_D6_reg  <= RDC1_D5_reg ;                   
 			RDC1_D7_reg  <= RDC1_D6_reg ;                   
 			RDC1_D8_reg  <= RDC1_D7_reg ;                   
 			RDC1_D9_reg  <= RDC1_D8_reg ;                   
 			RDC1_D10_reg <= RDC1_D9_reg ;                   
 			RDC1_D11_reg <= RDC1_D10_reg ;                  
 			RDC1_D12_reg <= RDC1_D11_reg ;                  
 			RDC1_D13_reg <= RDC1_D12_reg ;                  
 			RDC1_D14_reg <= RDC1_D13_reg ;                  
 			RDC1_D15_reg <= RDC1_D14_reg ;                  
 			RDC1_D16_reg <= RDC1_D15_reg ;                  
 			RDC1_D17_reg <= RDC1_D16_reg ;                  
 			RDC1_D18_reg <= RDC1_D17_reg ;                  
 			RDC1_D19_reg <= RDC1_D18_reg ;                  
 			RDC1_D20_reg <= RDC1_D19_reg ;                  
 			RDC1_D21_reg <= RDC1_D20_reg ;                  
 			RDC1_D_out   <= RDC1_D21_reg ;                  
 			//                                              
 			RDC2_D0_reg  <= RDC2_in ;                       
 			RDC2_D1_reg  <= RDC2_D0_reg ;                   
 			RDC2_D2_reg  <= RDC2_D1_reg ;                   
 			RDC2_D3_reg  <= RDC2_D2_reg ;                   
 			RDC2_D4_reg  <= RDC2_D3_reg ;                   
 			RDC2_D5_reg  <= RDC2_D4_reg ;                   
 			RDC2_D6_reg  <= RDC2_D5_reg ;                   
 			RDC2_D7_reg  <= RDC2_D6_reg ;                   
 			RDC2_D8_reg  <= RDC2_D7_reg ;                   
 			RDC2_D9_reg  <= RDC2_D8_reg ;                   
 			RDC2_D10_reg <= RDC2_D9_reg ;                   
 			RDC2_D11_reg <= RDC2_D10_reg ;                  
 			RDC2_D12_reg <= RDC2_D11_reg ;                  
 			RDC2_D13_reg <= RDC2_D12_reg ;                  
 			RDC2_D14_reg <= RDC2_D13_reg ;                  
 			RDC2_D15_reg <= RDC2_D14_reg ;                  
 			RDC2_D16_reg <= RDC2_D15_reg ;                  
 			RDC2_D17_reg <= RDC2_D16_reg ;                  
 			RDC2_D18_reg <= RDC2_D17_reg ;                  
 			RDC2_D19_reg <= RDC2_D18_reg ;                  
 			RDC2_D20_reg <= RDC2_D19_reg ;                  
 			RDC2_D21_reg <= RDC2_D20_reg ;                  
 			RDC2_D_out   <= RDC2_D21_reg ;                  
 			//                                              
 			RDC3_D0_reg  <= RDC3_in ;                       
 			RDC3_D1_reg  <= RDC3_D0_reg ;                   
 			RDC3_D2_reg  <= RDC3_D1_reg ;                   
 			RDC3_D3_reg  <= RDC3_D2_reg ;                   
 			RDC3_D4_reg  <= RDC3_D3_reg ;                   
 			RDC3_D5_reg  <= RDC3_D4_reg ;                   
 			RDC3_D6_reg  <= RDC3_D5_reg ;                   
 			RDC3_D7_reg  <= RDC3_D6_reg ;                   
 			RDC3_D8_reg  <= RDC3_D7_reg ;                   
 			RDC3_D9_reg  <= RDC3_D8_reg ;                   
 			RDC3_D10_reg <= RDC3_D9_reg ;                   
 			RDC3_D11_reg <= RDC3_D10_reg ;                  
 			RDC3_D12_reg <= RDC3_D11_reg ;                  
 			RDC3_D13_reg <= RDC3_D12_reg ;                  
 			RDC3_D14_reg <= RDC3_D13_reg ;                  
 			RDC3_D15_reg <= RDC3_D14_reg ;                  
 			RDC3_D16_reg <= RDC3_D15_reg ;                  
 			RDC3_D17_reg <= RDC3_D16_reg ;                  
 			RDC3_D18_reg <= RDC3_D17_reg ;                  
 			RDC3_D19_reg <= RDC3_D18_reg ;                  
 			RDC3_D20_reg <= RDC3_D19_reg ;                  
 			RDC3_D21_reg <= RDC3_D20_reg ;                  
 			RDC3_D_out   <= RDC3_D21_reg ;                  
 			//                                              
 			RDC4_D0_reg  <= RDC4_in ;                       
 			RDC4_D1_reg  <= RDC4_D0_reg ;                   
 			RDC4_D2_reg  <= RDC4_D1_reg ;                   
 			RDC4_D3_reg  <= RDC4_D2_reg ;                   
 			RDC4_D4_reg  <= RDC4_D3_reg ;                   
 			RDC4_D5_reg  <= RDC4_D4_reg ;                   
 			RDC4_D6_reg  <= RDC4_D5_reg ;                   
 			RDC4_D7_reg  <= RDC4_D6_reg ;                   
 			RDC4_D8_reg  <= RDC4_D7_reg ;                   
 			RDC4_D9_reg  <= RDC4_D8_reg ;                   
 			RDC4_D10_reg <= RDC4_D9_reg ;                   
 			RDC4_D11_reg <= RDC4_D10_reg ;                  
 			RDC4_D12_reg <= RDC4_D11_reg ;                  
 			RDC4_D13_reg <= RDC4_D12_reg ;                  
 			RDC4_D14_reg <= RDC4_D13_reg ;                  
 			RDC4_D15_reg <= RDC4_D14_reg ;                  
 			RDC4_D16_reg <= RDC4_D15_reg ;                  
 			RDC4_D17_reg <= RDC4_D16_reg ;                  
 			RDC4_D18_reg <= RDC4_D17_reg ;                  
 			RDC4_D19_reg <= RDC4_D18_reg ;                  
 			RDC4_D20_reg <= RDC4_D19_reg ;                  
 			RDC4_D21_reg <= RDC4_D20_reg ;                  
 			RDC4_D_out   <= RDC4_D21_reg ;                  
 			//                                              
 			RDC5_D0_reg  <= RDC5_in ;                       
 			RDC5_D1_reg  <= RDC5_D0_reg ;                   
 			RDC5_D2_reg  <= RDC5_D1_reg ;                   
 			RDC5_D3_reg  <= RDC5_D2_reg ;                   
 			RDC5_D4_reg  <= RDC5_D3_reg ;                   
 			RDC5_D5_reg  <= RDC5_D4_reg ;                   
 			RDC5_D6_reg  <= RDC5_D5_reg ;                   
 			RDC5_D7_reg  <= RDC5_D6_reg ;                   
 			RDC5_D8_reg  <= RDC5_D7_reg ;                   
 			RDC5_D9_reg  <= RDC5_D8_reg ;                   
 			RDC5_D10_reg <= RDC5_D9_reg ;                   
 			RDC5_D11_reg <= RDC5_D10_reg ;                  
 			RDC5_D12_reg <= RDC5_D11_reg ;                  
 			RDC5_D13_reg <= RDC5_D12_reg ;                  
 			RDC5_D14_reg <= RDC5_D13_reg ;                  
 			RDC5_D15_reg <= RDC5_D14_reg ;                  
 			RDC5_D16_reg <= RDC5_D15_reg ;                  
 			RDC5_D17_reg <= RDC5_D16_reg ;                  
 			RDC5_D18_reg <= RDC5_D17_reg ;                  
 			RDC5_D19_reg <= RDC5_D18_reg ;                  
 			RDC5_D20_reg <= RDC5_D19_reg ;                  
 			RDC5_D21_reg <= RDC5_D20_reg ;                  
 			RDC5_D_out   <= RDC5_D21_reg ;                  
 			//                                              
 			RDC6_D0_reg  <= RDC6_in ;                       
 			RDC6_D1_reg  <= RDC6_D0_reg ;                   
 			RDC6_D2_reg  <= RDC6_D1_reg ;                   
 			RDC6_D3_reg  <= RDC6_D2_reg ;                   
 			RDC6_D4_reg  <= RDC6_D3_reg ;                   
 			RDC6_D5_reg  <= RDC6_D4_reg ;                   
 			RDC6_D6_reg  <= RDC6_D5_reg ;                   
 			RDC6_D7_reg  <= RDC6_D6_reg ;                   
 			RDC6_D8_reg  <= RDC6_D7_reg ;                   
 			RDC6_D9_reg  <= RDC6_D8_reg ;                   
 			RDC6_D10_reg <= RDC6_D9_reg ;                   
 			RDC6_D11_reg <= RDC6_D10_reg ;                  
 			RDC6_D12_reg <= RDC6_D11_reg ;                  
 			RDC6_D13_reg <= RDC6_D12_reg ;                  
 			RDC6_D14_reg <= RDC6_D13_reg ;                  
 			RDC6_D15_reg <= RDC6_D14_reg ;                  
 			RDC6_D16_reg <= RDC6_D15_reg ;                  
 			RDC6_D17_reg <= RDC6_D16_reg ;                  
 			RDC6_D18_reg <= RDC6_D17_reg ;                  
 			RDC6_D19_reg <= RDC6_D18_reg ;                  
 			RDC6_D20_reg <= RDC6_D19_reg ;                  
 			RDC6_D21_reg <= RDC6_D20_reg ;                  
 			RDC6_D_out   <= RDC6_D21_reg ;                  
 			//                                              
 			RDC7_D0_reg  <= RDC7_in ;                       
 			RDC7_D1_reg  <= RDC7_D0_reg ;                   
 			RDC7_D2_reg  <= RDC7_D1_reg ;                   
 			RDC7_D3_reg  <= RDC7_D2_reg ;                   
 			RDC7_D4_reg  <= RDC7_D3_reg ;                   
 			RDC7_D5_reg  <= RDC7_D4_reg ;                   
 			RDC7_D6_reg  <= RDC7_D5_reg ;                   
 			RDC7_D7_reg  <= RDC7_D6_reg ;                   
 			RDC7_D8_reg  <= RDC7_D7_reg ;                   
 			RDC7_D9_reg  <= RDC7_D8_reg ;                   
 			RDC7_D10_reg <= RDC7_D9_reg ;                   
 			RDC7_D11_reg <= RDC7_D10_reg ;                  
 			RDC7_D12_reg <= RDC7_D11_reg ;                  
 			RDC7_D13_reg <= RDC7_D12_reg ;                  
 			RDC7_D14_reg <= RDC7_D13_reg ;                  
 			RDC7_D15_reg <= RDC7_D14_reg ;                  
 			RDC7_D16_reg <= RDC7_D15_reg ;                  
 			RDC7_D17_reg <= RDC7_D16_reg ;                  
 			RDC7_D18_reg <= RDC7_D17_reg ;                  
 			RDC7_D19_reg <= RDC7_D18_reg ;                  
 			RDC7_D20_reg <= RDC7_D19_reg ;                  
 			RDC7_D21_reg <= RDC7_D20_reg ;                  
 			RDC7_D_out   <= RDC7_D21_reg ;                  
 			//                                              
 			RDC8_D0_reg  <= RDC8_in ;                       
 			RDC8_D1_reg  <= RDC8_D0_reg ;                   
 			RDC8_D2_reg  <= RDC8_D1_reg ;                   
 			RDC8_D3_reg  <= RDC8_D2_reg ;                   
 			RDC8_D4_reg  <= RDC8_D3_reg ;                   
 			RDC8_D5_reg  <= RDC8_D4_reg ;                   
 			RDC8_D6_reg  <= RDC8_D5_reg ;                   
 			RDC8_D7_reg  <= RDC8_D6_reg ;                   
 			RDC8_D8_reg  <= RDC8_D7_reg ;                   
 			RDC8_D9_reg  <= RDC8_D8_reg ;                   
 			RDC8_D10_reg <= RDC8_D9_reg ;                   
 			RDC8_D11_reg <= RDC8_D10_reg ;                  
 			RDC8_D12_reg <= RDC8_D11_reg ;                  
 			RDC8_D13_reg <= RDC8_D12_reg ;                  
 			RDC8_D14_reg <= RDC8_D13_reg ;                  
 			RDC8_D15_reg <= RDC8_D14_reg ;                  
 			RDC8_D16_reg <= RDC8_D15_reg ;                  
 			RDC8_D17_reg <= RDC8_D16_reg ;                  
 			RDC8_D18_reg <= RDC8_D17_reg ;                  
 			RDC8_D19_reg <= RDC8_D18_reg ;                  
 			RDC8_D20_reg <= RDC8_D19_reg ;                  
 			RDC8_D21_reg <= RDC8_D20_reg ;                  
 			RDC8_D_out   <= RDC8_D21_reg ;                  
 			//                                              
 			RDC9_D0_reg  <= RDC9_in ;                       
 			RDC9_D1_reg  <= RDC9_D0_reg ;                   
 			RDC9_D2_reg  <= RDC9_D1_reg ;                   
 			RDC9_D3_reg  <= RDC9_D2_reg ;                   
 			RDC9_D4_reg  <= RDC9_D3_reg ;                   
 			RDC9_D5_reg  <= RDC9_D4_reg ;                   
 			RDC9_D6_reg  <= RDC9_D5_reg ;                   
 			RDC9_D7_reg  <= RDC9_D6_reg ;                   
 			RDC9_D8_reg  <= RDC9_D7_reg ;                   
 			RDC9_D9_reg  <= RDC9_D8_reg ;                   
 			RDC9_D10_reg <= RDC9_D9_reg ;                   
 			RDC9_D11_reg <= RDC9_D10_reg ;                  
 			RDC9_D12_reg <= RDC9_D11_reg ;                  
 			RDC9_D13_reg <= RDC9_D12_reg ;                  
 			RDC9_D14_reg <= RDC9_D13_reg ;                  
 			RDC9_D15_reg <= RDC9_D14_reg ;                  
 			RDC9_D16_reg <= RDC9_D15_reg ;                  
 			RDC9_D17_reg <= RDC9_D16_reg ;                  
 			RDC9_D18_reg <= RDC9_D17_reg ;                  
 			RDC9_D19_reg <= RDC9_D18_reg ;                  
 			RDC9_D20_reg <= RDC9_D19_reg ;                  
 			RDC9_D21_reg <= RDC9_D20_reg ;                  
 			RDC9_D_out   <= RDC9_D21_reg ;                  
 			//                                              
 			RDC10_D0_reg  <= RDC10_in ;                     
 			RDC10_D1_reg  <= RDC10_D0_reg ;                 
 			RDC10_D2_reg  <= RDC10_D1_reg ;                 
 			RDC10_D3_reg  <= RDC10_D2_reg ;                 
 			RDC10_D4_reg  <= RDC10_D3_reg ;                 
 			RDC10_D5_reg  <= RDC10_D4_reg ;                 
 			RDC10_D6_reg  <= RDC10_D5_reg ;                 
 			RDC10_D7_reg  <= RDC10_D6_reg ;                 
 			RDC10_D8_reg  <= RDC10_D7_reg ;                 
 			RDC10_D9_reg  <= RDC10_D8_reg ;                 
 			RDC10_D10_reg <= RDC10_D9_reg ;                 
 			RDC10_D11_reg <= RDC10_D10_reg ;                
 			RDC10_D12_reg <= RDC10_D11_reg ;                
 			RDC10_D13_reg <= RDC10_D12_reg ;                
 			RDC10_D14_reg <= RDC10_D13_reg ;                
 			RDC10_D15_reg <= RDC10_D14_reg ;                
 			RDC10_D16_reg <= RDC10_D15_reg ;                
 			RDC10_D17_reg <= RDC10_D16_reg ;                
 			RDC10_D18_reg <= RDC10_D17_reg ;                
 			RDC10_D19_reg <= RDC10_D18_reg ;                
 			RDC10_D20_reg <= RDC10_D19_reg ;                
 			RDC10_D21_reg <= RDC10_D20_reg ;                
 			RDC10_D_out   <= RDC10_D21_reg ;                
 			//                                              
 			RDC11_D0_reg  <= RDC11_in ;                     
 			RDC11_D1_reg  <= RDC11_D0_reg ;                 
 			RDC11_D2_reg  <= RDC11_D1_reg ;                 
 			RDC11_D3_reg  <= RDC11_D2_reg ;                 
 			RDC11_D4_reg  <= RDC11_D3_reg ;                 
 			RDC11_D5_reg  <= RDC11_D4_reg ;                 
 			RDC11_D6_reg  <= RDC11_D5_reg ;                 
 			RDC11_D7_reg  <= RDC11_D6_reg ;                 
 			RDC11_D8_reg  <= RDC11_D7_reg ;                 
 			RDC11_D9_reg  <= RDC11_D8_reg ;                 
 			RDC11_D10_reg <= RDC11_D9_reg ;                 
 			RDC11_D11_reg <= RDC11_D10_reg ;                
 			RDC11_D12_reg <= RDC11_D11_reg ;                
 			RDC11_D13_reg <= RDC11_D12_reg ;                
 			RDC11_D14_reg <= RDC11_D13_reg ;                
 			RDC11_D15_reg <= RDC11_D14_reg ;                
 			RDC11_D16_reg <= RDC11_D15_reg ;                
 			RDC11_D17_reg <= RDC11_D16_reg ;                
 			RDC11_D18_reg <= RDC11_D17_reg ;                
 			RDC11_D19_reg <= RDC11_D18_reg ;                
 			RDC11_D20_reg <= RDC11_D19_reg ;                
 			RDC11_D21_reg <= RDC11_D20_reg ;                
 			RDC11_D_out   <= RDC11_D21_reg ;                
 			//                                              
 			RDC12_D0_reg  <= RDC12_in ;                     
 			RDC12_D1_reg  <= RDC12_D0_reg ;                 
 			RDC12_D2_reg  <= RDC12_D1_reg ;                 
 			RDC12_D3_reg  <= RDC12_D2_reg ;                 
 			RDC12_D4_reg  <= RDC12_D3_reg ;                 
 			RDC12_D5_reg  <= RDC12_D4_reg ;                 
 			RDC12_D6_reg  <= RDC12_D5_reg ;                 
 			RDC12_D7_reg  <= RDC12_D6_reg ;                 
 			RDC12_D8_reg  <= RDC12_D7_reg ;                 
 			RDC12_D9_reg  <= RDC12_D8_reg ;                 
 			RDC12_D10_reg <= RDC12_D9_reg ;                 
 			RDC12_D11_reg <= RDC12_D10_reg ;                
 			RDC12_D12_reg <= RDC12_D11_reg ;                
 			RDC12_D13_reg <= RDC12_D12_reg ;                
 			RDC12_D14_reg <= RDC12_D13_reg ;                
 			RDC12_D15_reg <= RDC12_D14_reg ;                
 			RDC12_D16_reg <= RDC12_D15_reg ;                
 			RDC12_D17_reg <= RDC12_D16_reg ;                
 			RDC12_D18_reg <= RDC12_D17_reg ;                
 			RDC12_D19_reg <= RDC12_D18_reg ;                
 			RDC12_D20_reg <= RDC12_D19_reg ;                
 			RDC12_D21_reg <= RDC12_D20_reg ;                
 			RDC12_D_out   <= RDC12_D21_reg ;                
 			//                                              
 			RDC13_D0_reg  <= RDC13_in ;                     
 			RDC13_D1_reg  <= RDC13_D0_reg ;                 
 			RDC13_D2_reg  <= RDC13_D1_reg ;                 
 			RDC13_D3_reg  <= RDC13_D2_reg ;                 
 			RDC13_D4_reg  <= RDC13_D3_reg ;                 
 			RDC13_D5_reg  <= RDC13_D4_reg ;                 
 			RDC13_D6_reg  <= RDC13_D5_reg ;                 
 			RDC13_D7_reg  <= RDC13_D6_reg ;                 
 			RDC13_D8_reg  <= RDC13_D7_reg ;                 
 			RDC13_D9_reg  <= RDC13_D8_reg ;                 
 			RDC13_D10_reg <= RDC13_D9_reg ;                 
 			RDC13_D11_reg <= RDC13_D10_reg ;                
 			RDC13_D12_reg <= RDC13_D11_reg ;                
 			RDC13_D13_reg <= RDC13_D12_reg ;                
 			RDC13_D14_reg <= RDC13_D13_reg ;                
 			RDC13_D15_reg <= RDC13_D14_reg ;                
 			RDC13_D16_reg <= RDC13_D15_reg ;                
 			RDC13_D17_reg <= RDC13_D16_reg ;                
 			RDC13_D18_reg <= RDC13_D17_reg ;                
 			RDC13_D19_reg <= RDC13_D18_reg ;                
 			RDC13_D20_reg <= RDC13_D19_reg ;                
 			RDC13_D21_reg <= RDC13_D20_reg ;                
 			RDC13_D_out   <= RDC13_D21_reg ;                
 			//                                              
 			RDC14_D0_reg  <= RDC14_in ;                     
 			RDC14_D1_reg  <= RDC14_D0_reg ;                 
 			RDC14_D2_reg  <= RDC14_D1_reg ;                 
 			RDC14_D3_reg  <= RDC14_D2_reg ;                 
 			RDC14_D4_reg  <= RDC14_D3_reg ;                 
 			RDC14_D5_reg  <= RDC14_D4_reg ;                 
 			RDC14_D6_reg  <= RDC14_D5_reg ;                 
 			RDC14_D7_reg  <= RDC14_D6_reg ;                 
 			RDC14_D8_reg  <= RDC14_D7_reg ;                 
 			RDC14_D9_reg  <= RDC14_D8_reg ;                 
 			RDC14_D10_reg <= RDC14_D9_reg ;                 
 			RDC14_D11_reg <= RDC14_D10_reg ;                
 			RDC14_D12_reg <= RDC14_D11_reg ;                
 			RDC14_D13_reg <= RDC14_D12_reg ;                
 			RDC14_D14_reg <= RDC14_D13_reg ;                
 			RDC14_D15_reg <= RDC14_D14_reg ;                
 			RDC14_D16_reg <= RDC14_D15_reg ;                
 			RDC14_D17_reg <= RDC14_D16_reg ;                
 			RDC14_D18_reg <= RDC14_D17_reg ;                
 			RDC14_D19_reg <= RDC14_D18_reg ;                
 			RDC14_D20_reg <= RDC14_D19_reg ;                
 			RDC14_D21_reg <= RDC14_D20_reg ;                
 			RDC14_D_out   <= RDC14_D21_reg ;                
 			//                                              
 			RDC15_D0_reg  <= RDC15_in ;                     
 			RDC15_D1_reg  <= RDC15_D0_reg ;                 
 			RDC15_D2_reg  <= RDC15_D1_reg ;                 
 			RDC15_D3_reg  <= RDC15_D2_reg ;                 
 			RDC15_D4_reg  <= RDC15_D3_reg ;                 
 			RDC15_D5_reg  <= RDC15_D4_reg ;                 
 			RDC15_D6_reg  <= RDC15_D5_reg ;                 
 			RDC15_D7_reg  <= RDC15_D6_reg ;                 
 			RDC15_D8_reg  <= RDC15_D7_reg ;                 
 			RDC15_D9_reg  <= RDC15_D8_reg ;                 
 			RDC15_D10_reg <= RDC15_D9_reg ;                 
 			RDC15_D11_reg <= RDC15_D10_reg ;                
 			RDC15_D12_reg <= RDC15_D11_reg ;                
 			RDC15_D13_reg <= RDC15_D12_reg ;                
 			RDC15_D14_reg <= RDC15_D13_reg ;                
 			RDC15_D15_reg <= RDC15_D14_reg ;                
 			RDC15_D16_reg <= RDC15_D15_reg ;                
 			RDC15_D17_reg <= RDC15_D16_reg ;                
 			RDC15_D18_reg <= RDC15_D17_reg ;                
 			RDC15_D19_reg <= RDC15_D18_reg ;                
 			RDC15_D20_reg <= RDC15_D19_reg ;                
 			RDC15_D21_reg <= RDC15_D20_reg ;                
 			RDC15_D_out   <= RDC15_D21_reg ;                
 		end                                                 
 	end                                                     
 endmodule                                                   
