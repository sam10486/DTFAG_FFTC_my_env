`include "define.v"
module Memory_wrapper (
    input clk,
    input rst_n,
    input ROM_CEN,
    input [1:0] FFT_stage_in,
    input [`ROMA_width-1:0] MA0,
    input [`ROMA_width-1:0] MA1,
    input [`ROMA_width-1:0] MA2,

    output wire [`D_width-1:0] ROM0_b0   ,
    output wire [`D_width-1:0] ROM0_b1   ,
    output wire [`D_width-1:0] ROM0_b2   ,
    output wire [`D_width-1:0] ROM0_b3   ,
    output wire [`D_width-1:0] ROM0_b4   ,
    output wire [`D_width-1:0] ROM0_b5   ,
    output wire [`D_width-1:0] ROM0_b6   ,
    output wire [`D_width-1:0] ROM0_b7   ,
    output wire [`D_width-1:0] ROM0_b8   ,
    output wire [`D_width-1:0] ROM0_b9   ,
    output wire [`D_width-1:0] ROM0_b10  ,
    output wire [`D_width-1:0] ROM0_b11  ,
    output wire [`D_width-1:0] ROM0_b12  ,
    output wire [`D_width-1:0] ROM0_b13  ,
    output wire [`D_width-1:0] ROM0_b14  ,
    output wire [`D_width-1:0] ROM0_b15  ,
    // ROM1
    output wire [`D_width-1:0] ROM1_b0   ,
    output wire [`D_width-1:0] ROM1_b1   ,
    output wire [`D_width-1:0] ROM1_b2   ,
    output wire [`D_width-1:0] ROM1_b3   ,
    output wire [`D_width-1:0] ROM1_b4   ,
    output wire [`D_width-1:0] ROM1_b5   ,
    output wire [`D_width-1:0] ROM1_b6   ,
    output wire [`D_width-1:0] ROM1_b7   ,
    output wire [`D_width-1:0] ROM1_b8   ,
    output wire [`D_width-1:0] ROM1_b9   ,
    output wire [`D_width-1:0] ROM1_b10  ,
    output wire [`D_width-1:0] ROM1_b11  ,
    output wire [`D_width-1:0] ROM1_b12  ,
    output wire [`D_width-1:0] ROM1_b13  ,
    output wire [`D_width-1:0] ROM1_b14  ,
    output wire [`D_width-1:0] ROM1_b15  ,
    // ROM2
    output wire [`D_width-1:0] ROM2_b0   ,
    output wire [`D_width-1:0] ROM2_b1   ,
    output wire [`D_width-1:0] ROM2_b2   ,
    output wire [`D_width-1:0] ROM2_b3   ,
    output wire [`D_width-1:0] ROM2_b4   ,
    output wire [`D_width-1:0] ROM2_b5   ,
    output wire [`D_width-1:0] ROM2_b6   ,
    output wire [`D_width-1:0] ROM2_b7   ,
    output wire [`D_width-1:0] ROM2_b8   ,
    output wire [`D_width-1:0] ROM2_b9   ,
    output wire [`D_width-1:0] ROM2_b10  ,
    output wire [`D_width-1:0] ROM2_b11  ,
    output wire [`D_width-1:0] ROM2_b12  ,
    output wire [`D_width-1:0] ROM2_b13  ,
    output wire [`D_width-1:0] ROM2_b14  ,
    output wire [`D_width-1:0] ROM2_b15  

);

    
    Register_file Register_file(
        .clk       (clk     ),
        .rst_n     (rst_n   ),
        .MA0       (MA0     ),
        .MA1       (MA1     ),
        .MA2       (MA2     ),
        .ROM_CEN   (ROM_CEN ),
        .FFT_stage_in(FFT_stage_in),
        // output
        // ROM0
        .ROM0_b0   (ROM0_b0 ),
        .ROM0_b1   (ROM0_b1 ),
        .ROM0_b2   (ROM0_b2 ),
        .ROM0_b3   (ROM0_b3 ),
        .ROM0_b4   (ROM0_b4 ),
        .ROM0_b5   (ROM0_b5 ),
        .ROM0_b6   (ROM0_b6 ),
        .ROM0_b7   (ROM0_b7 ),
        .ROM0_b8   (ROM0_b8 ),
        .ROM0_b9   (ROM0_b9 ),
        .ROM0_b10  (ROM0_b10),
        .ROM0_b11  (ROM0_b11),
        .ROM0_b12  (ROM0_b12),
        .ROM0_b13  (ROM0_b13),
        .ROM0_b14  (ROM0_b14),
        .ROM0_b15  (ROM0_b15),
        // ROM1
        .ROM1_b0   (ROM1_b0 ),
        .ROM1_b1   (ROM1_b1 ),
        .ROM1_b2   (ROM1_b2 ),
        .ROM1_b3   (ROM1_b3 ),
        .ROM1_b4   (ROM1_b4 ),
        .ROM1_b5   (ROM1_b5 ),
        .ROM1_b6   (ROM1_b6 ),
        .ROM1_b7   (ROM1_b7 ),
        .ROM1_b8   (ROM1_b8 ),
        .ROM1_b9   (ROM1_b9 ),
        .ROM1_b10  (ROM1_b10),
        .ROM1_b11  (ROM1_b11),
        .ROM1_b12  (ROM1_b12),
        .ROM1_b13  (ROM1_b13),
        .ROM1_b14  (ROM1_b14),
        .ROM1_b15  (ROM1_b15),
        // ROM2
        .ROM2_b0   (ROM2_b0 ),
        .ROM2_b1   (ROM2_b1 ),
        .ROM2_b2   (ROM2_b2 ),
        .ROM2_b3   (ROM2_b3 ),
        .ROM2_b4   (ROM2_b4 ),
        .ROM2_b5   (ROM2_b5 ),
        .ROM2_b6   (ROM2_b6 ),
        .ROM2_b7   (ROM2_b7 ),
        .ROM2_b8   (ROM2_b8 ),
        .ROM2_b9   (ROM2_b9 ),
        .ROM2_b10  (ROM2_b10),
        .ROM2_b11  (ROM2_b11),
        .ROM2_b12  (ROM2_b12),
        .ROM2_b13  (ROM2_b13),
        .ROM2_b14  (ROM2_b14),
        .ROM2_b15  (ROM2_b15)
    );



endmodule