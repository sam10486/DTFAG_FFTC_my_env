`include "define.v"
module Register_file (
    input clk,
    input rst_n,
    input [`ROMA_width-1:0] MA0,
    input [`ROMA_width-1:0] MA1,
    input [`ROMA_width-1:0] MA2,
    input ROM_CEN,

    output reg [`D_width-1:0] ROM0_b0   ,
    output reg [`D_width-1:0] ROM0_b1   ,
    output reg [`D_width-1:0] ROM0_b2   ,
    output reg [`D_width-1:0] ROM0_b3   ,
    output reg [`D_width-1:0] ROM0_b4   ,
    output reg [`D_width-1:0] ROM0_b5   ,
    output reg [`D_width-1:0] ROM0_b6   ,
    output reg [`D_width-1:0] ROM0_b7   ,
    output reg [`D_width-1:0] ROM0_b8   ,
    output reg [`D_width-1:0] ROM0_b9   ,
    output reg [`D_width-1:0] ROM0_b10  ,
    output reg [`D_width-1:0] ROM0_b11  ,
    output reg [`D_width-1:0] ROM0_b12  ,
    output reg [`D_width-1:0] ROM0_b13  ,
    output reg [`D_width-1:0] ROM0_b14  ,
    output reg [`D_width-1:0] ROM0_b15  ,
    // ROM1
    output reg [`D_width-1:0] ROM1_b0   ,
    output reg [`D_width-1:0] ROM1_b1   ,
    output reg [`D_width-1:0] ROM1_b2   ,
    output reg [`D_width-1:0] ROM1_b3   ,
    output reg [`D_width-1:0] ROM1_b4   ,
    output reg [`D_width-1:0] ROM1_b5   ,
    output reg [`D_width-1:0] ROM1_b6   ,
    output reg [`D_width-1:0] ROM1_b7   ,
    output reg [`D_width-1:0] ROM1_b8   ,
    output reg [`D_width-1:0] ROM1_b9   ,
    output reg [`D_width-1:0] ROM1_b10  ,
    output reg [`D_width-1:0] ROM1_b11  ,
    output reg [`D_width-1:0] ROM1_b12  ,
    output reg [`D_width-1:0] ROM1_b13  ,
    output reg [`D_width-1:0] ROM1_b14  ,
    output reg [`D_width-1:0] ROM1_b15  ,
    // ROM2
    output reg [`D_width-1:0] ROM2_b0   ,
    output reg [`D_width-1:0] ROM2_b1   ,
    output reg [`D_width-1:0] ROM2_b2   ,
    output reg [`D_width-1:0] ROM2_b3   ,
    output reg [`D_width-1:0] ROM2_b4   ,
    output reg [`D_width-1:0] ROM2_b5   ,
    output reg [`D_width-1:0] ROM2_b6   ,
    output reg [`D_width-1:0] ROM2_b7   ,
    output reg [`D_width-1:0] ROM2_b8   ,
    output reg [`D_width-1:0] ROM2_b9   ,
    output reg [`D_width-1:0] ROM2_b10  ,
    output reg [`D_width-1:0] ROM2_b11  ,
    output reg [`D_width-1:0] ROM2_b12  ,
    output reg [`D_width-1:0] ROM2_b13  ,
    output reg [`D_width-1:0] ROM2_b14  ,
    output reg [`D_width-1:0] ROM2_b15  
);

    reg [`D_width-1:0] ROM0_arr [0:15][0:15];
    reg [`D_width-1:0] ROM1_arr [0:15][0:15];
    reg [`D_width-1:0] ROM2_arr [0:15][0:15];
    
    always@( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            // ROM0 init
            ROM0_arr[0][0] <= 64'd1;
            ROM0_arr[1][0] <= 64'd1;
            ROM0_arr[2][0] <= 64'd1;
            ROM0_arr[3][0] <= 64'd1;
            ROM0_arr[4][0] <= 64'd1;
            ROM0_arr[5][0] <= 64'd1;
            ROM0_arr[6][0] <= 64'd1;
            ROM0_arr[7][0] <= 64'd1;
            ROM0_arr[8][0] <= 64'd1;
            ROM0_arr[9][0] <= 64'd1;
            ROM0_arr[10][0] <= 64'd1;
            ROM0_arr[11][0] <= 64'd1;
            ROM0_arr[12][0] <= 64'd1;
            ROM0_arr[13][0] <= 64'd1;
            ROM0_arr[14][0] <= 64'd1;
            ROM0_arr[15][0] <= 64'd1;
            ROM0_arr[0][1] <= 64'd1;
            ROM0_arr[1][1] <= 64'd11147770252432840497;
            ROM0_arr[2][1] <= 64'd18446181119461163011;
            ROM0_arr[3][1] <= 64'd6562114217670983589;
            ROM0_arr[4][1] <= 64'd18444492269600899073;
            ROM0_arr[5][1] <= 64'd10853271128879547664;
            ROM0_arr[6][1] <= 64'd18442240469787213809;
            ROM0_arr[7][1] <= 64'd9362914843564906265;
            ROM0_arr[8][1] <= 64'd18446744069414584257;
            ROM0_arr[9][1] <= 64'd5965722551466996711;
            ROM0_arr[10][1] <= 64'd36028797018963840;
            ROM0_arr[11][1] <= 64'd4299803665592489687;
            ROM0_arr[12][1] <= 64'd144115188075855872;
            ROM0_arr[13][1] <= 64'd6366922389463153702;
            ROM0_arr[14][1] <= 64'd288230376151712768;
            ROM0_arr[15][1] <= 64'd9516004302527281633;
            ROM0_arr[0][2] <= 64'd1;
            ROM0_arr[1][2] <= 64'd18446181119461163011;
            ROM0_arr[2][2] <= 64'd18444492269600899073;
            ROM0_arr[3][2] <= 64'd18442240469787213809;
            ROM0_arr[4][2] <= 64'd18446744069414584257;
            ROM0_arr[5][2] <= 64'd36028797018963840;
            ROM0_arr[6][2] <= 64'd144115188075855872;
            ROM0_arr[7][2] <= 64'd288230376151712768;
            ROM0_arr[8][2] <= 64'd4096;
            ROM0_arr[9][2] <= 64'd16140901060200898561;
            ROM0_arr[10][2] <= 64'd9223372032559808513;
            ROM0_arr[11][2] <= 64'd18446744065119551490;
            ROM0_arr[12][2] <= 64'd18446744069414322177;
            ROM0_arr[13][2] <= 64'd34359214072;
            ROM0_arr[14][2] <= 64'd137438953440;
            ROM0_arr[15][2] <= 64'd274882101184;
            ROM0_arr[0][3] <= 64'd1;
            ROM0_arr[1][3] <= 64'd6562114217670983589;
            ROM0_arr[2][3] <= 64'd18442240469787213809;
            ROM0_arr[3][3] <= 64'd5965722551466996711;
            ROM0_arr[4][3] <= 64'd144115188075855872;
            ROM0_arr[5][3] <= 64'd9516004302527281633;
            ROM0_arr[6][3] <= 64'd16140901060200898561;
            ROM0_arr[7][3] <= 64'd16792080670893602455;
            ROM0_arr[8][3] <= 64'd18446744069414322177;
            ROM0_arr[9][3] <= 64'd13801972045324315718;
            ROM0_arr[10][3] <= 64'd274882101184;
            ROM0_arr[11][3] <= 64'd18142929134658341675;
            ROM0_arr[12][3] <= 64'd18446735273321564161;
            ROM0_arr[13][3] <= 64'd8215369291935911999;
            ROM0_arr[14][3] <= 64'd140735340838912;
            ROM0_arr[15][3] <= 64'd3341893669734556710;
            ROM0_arr[0][4] <= 64'd1;
            ROM0_arr[1][4] <= 64'd18444492269600899073;
            ROM0_arr[2][4] <= 64'd18446744069414584257;
            ROM0_arr[3][4] <= 64'd144115188075855872;
            ROM0_arr[4][4] <= 64'd4096;
            ROM0_arr[5][4] <= 64'd9223372032559808513;
            ROM0_arr[6][4] <= 64'd18446744069414322177;
            ROM0_arr[7][4] <= 64'd137438953440;
            ROM0_arr[8][4] <= 64'd16777216;
            ROM0_arr[9][4] <= 64'd18446735273321564161;
            ROM0_arr[10][4] <= 64'd18446744068340842497;
            ROM0_arr[11][4] <= 64'd562949953290240;
            ROM0_arr[12][4] <= 64'd68719476736;
            ROM0_arr[13][4] <= 64'd18410715272404008961;
            ROM0_arr[14][4] <= 64'd18446739671368073217;
            ROM0_arr[15][4] <= 64'd2305843008676823040;
            ROM0_arr[0][5] <= 64'd1;
            ROM0_arr[1][5] <= 64'd10853271128879547664;
            ROM0_arr[2][5] <= 64'd36028797018963840;
            ROM0_arr[3][5] <= 64'd9516004302527281633;
            ROM0_arr[4][5] <= 64'd9223372032559808513;
            ROM0_arr[5][5] <= 64'd12110422903908887252;
            ROM0_arr[6][5] <= 64'd274882101184;
            ROM0_arr[7][5] <= 64'd2117504431143841456;
            ROM0_arr[8][5] <= 64'd18446744068340842497;
            ROM0_arr[9][5] <= 64'd3341893669734556710;
            ROM0_arr[10][5] <= 64'd18437737007600893953;
            ROM0_arr[11][5] <= 64'd3291437157293746400;
            ROM0_arr[12][5] <= 64'd2305843008676823040;
            ROM0_arr[13][5] <= 64'd17090085178304640863;
            ROM0_arr[14][5] <= 64'd18442240469787213841;
            ROM0_arr[15][5] <= 64'd1116342470860912836;
            ROM0_arr[0][6] <= 64'd1;
            ROM0_arr[1][6] <= 64'd18442240469787213809;
            ROM0_arr[2][6] <= 64'd144115188075855872;
            ROM0_arr[3][6] <= 64'd16140901060200898561;
            ROM0_arr[4][6] <= 64'd18446744069414322177;
            ROM0_arr[5][6] <= 64'd274882101184;
            ROM0_arr[6][6] <= 64'd18446735273321564161;
            ROM0_arr[7][6] <= 64'd140735340838912;
            ROM0_arr[8][6] <= 64'd68719476736;
            ROM0_arr[9][6] <= 64'd18374685375881805825;
            ROM0_arr[10][6] <= 64'd2305843008676823040;
            ROM0_arr[11][6] <= 64'd562949953421314;
            ROM0_arr[12][6] <= 64'd18428729670905102337;
            ROM0_arr[13][6] <= 64'd288230376151710720;
            ROM0_arr[14][6] <= 64'd32768;
            ROM0_arr[15][6] <= 64'd18446744035054321673;
            ROM0_arr[0][7] <= 64'd1;
            ROM0_arr[1][7] <= 64'd9362914843564906265;
            ROM0_arr[2][7] <= 64'd288230376151712768;
            ROM0_arr[3][7] <= 64'd16792080670893602455;
            ROM0_arr[4][7] <= 64'd137438953440;
            ROM0_arr[5][7] <= 64'd2117504431143841456;
            ROM0_arr[6][7] <= 64'd140735340838912;
            ROM0_arr[7][7] <= 64'd9952623958621855812;
            ROM0_arr[8][7] <= 64'd18446739671368073217;
            ROM0_arr[9][7] <= 64'd10708950766175242252;
            ROM0_arr[10][7] <= 64'd18442240469787213841;
            ROM0_arr[11][7] <= 64'd10832292272906805046;
            ROM0_arr[12][7] <= 64'd32768;
            ROM0_arr[13][7] <= 64'd16192975500896648969;
            ROM0_arr[14][7] <= 64'd2199056809472;
            ROM0_arr[15][7] <= 64'd13417321343344118652;
            ROM0_arr[0][8] <= 64'd1;
            ROM0_arr[1][8] <= 64'd18446744069414584257;
            ROM0_arr[2][8] <= 64'd4096;
            ROM0_arr[3][8] <= 64'd18446744069414322177;
            ROM0_arr[4][8] <= 64'd16777216;
            ROM0_arr[5][8] <= 64'd18446744068340842497;
            ROM0_arr[6][8] <= 64'd68719476736;
            ROM0_arr[7][8] <= 64'd18446739671368073217;
            ROM0_arr[8][8] <= 64'd281474976710656;
            ROM0_arr[9][8] <= 64'd18428729670905102337;
            ROM0_arr[10][8] <= 64'd1152921504606846976;
            ROM0_arr[11][8] <= 64'd18446744052234715141;
            ROM0_arr[12][8] <= 64'd1099511627520;
            ROM0_arr[13][8] <= 64'd18446673700670423041;
            ROM0_arr[14][8] <= 64'd4503599626321920;
            ROM0_arr[15][8] <= 64'd18158513693329981441;
            ROM0_arr[0][9] <= 64'd1;
            ROM0_arr[1][9] <= 64'd5965722551466996711;
            ROM0_arr[2][9] <= 64'd16140901060200898561;
            ROM0_arr[3][9] <= 64'd13801972045324315718;
            ROM0_arr[4][9] <= 64'd18446735273321564161;
            ROM0_arr[5][9] <= 64'd3341893669734556710;
            ROM0_arr[6][9] <= 64'd18374685375881805825;
            ROM0_arr[7][9] <= 64'd10708950766175242252;
            ROM0_arr[8][9] <= 64'd18428729670905102337;
            ROM0_arr[9][9] <= 64'd14041890976876060974;
            ROM0_arr[10][9] <= 64'd18446744035054321673;
            ROM0_arr[11][9] <= 64'd15113979899245772281;
            ROM0_arr[12][9] <= 64'd18446744060824649729;
            ROM0_arr[13][9] <= 64'd5834015391316509212;
            ROM0_arr[14][9] <= 64'd4611615648609468416;
            ROM0_arr[15][9] <= 64'd9083829225849678056;
            ROM0_arr[0][10] <= 64'd1;
            ROM0_arr[1][10] <= 64'd36028797018963840;
            ROM0_arr[2][10] <= 64'd9223372032559808513;
            ROM0_arr[3][10] <= 64'd274882101184;
            ROM0_arr[4][10] <= 64'd18446744068340842497;
            ROM0_arr[5][10] <= 64'd18437737007600893953;
            ROM0_arr[6][10] <= 64'd2305843008676823040;
            ROM0_arr[7][10] <= 64'd18442240469787213841;
            ROM0_arr[8][10] <= 64'd1152921504606846976;
            ROM0_arr[9][10] <= 64'd18446744035054321673;
            ROM0_arr[10][10] <= 64'd134217728;
            ROM0_arr[11][10] <= 64'd1125882726711296;
            ROM0_arr[12][10] <= 64'd18158513693329981441;
            ROM0_arr[13][10] <= 64'd562949953421310;
            ROM0_arr[14][10] <= 64'd18302628881338728449;
            ROM0_arr[15][10] <= 64'd4295032831;
            ROM0_arr[0][11] <= 64'd1;
            ROM0_arr[1][11] <= 64'd4299803665592489687;
            ROM0_arr[2][11] <= 64'd18446744065119551490;
            ROM0_arr[3][11] <= 64'd18142929134658341675;
            ROM0_arr[4][11] <= 64'd562949953290240;
            ROM0_arr[5][11] <= 64'd3291437157293746400;
            ROM0_arr[6][11] <= 64'd562949953421314;
            ROM0_arr[7][11] <= 64'd10832292272906805046;
            ROM0_arr[8][11] <= 64'd18446744052234715141;
            ROM0_arr[9][11] <= 64'd15113979899245772281;
            ROM0_arr[10][11] <= 64'd1125882726711296;
            ROM0_arr[11][11] <= 64'd4497639551463306333;
            ROM0_arr[12][11] <= 64'd2251799813685248;
            ROM0_arr[13][11] <= 64'd8930739766887302688;
            ROM0_arr[14][11] <= 64'd18446744035055370249;
            ROM0_arr[15][11] <= 64'd7546206866789277329;
            ROM0_arr[0][12] <= 64'd1;
            ROM0_arr[1][12] <= 64'd144115188075855872;
            ROM0_arr[2][12] <= 64'd18446744069414322177;
            ROM0_arr[3][12] <= 64'd18446735273321564161;
            ROM0_arr[4][12] <= 64'd68719476736;
            ROM0_arr[5][12] <= 64'd2305843008676823040;
            ROM0_arr[6][12] <= 64'd18428729670905102337;
            ROM0_arr[7][12] <= 64'd32768;
            ROM0_arr[8][12] <= 64'd1099511627520;
            ROM0_arr[9][12] <= 64'd18446744060824649729;
            ROM0_arr[10][12] <= 64'd18158513693329981441;
            ROM0_arr[11][12] <= 64'd2251799813685248;
            ROM0_arr[12][12] <= 64'd18446744069414580225;
            ROM0_arr[13][12] <= 64'd18446743931975630881;
            ROM0_arr[14][12] <= 64'd1073741824;
            ROM0_arr[15][12] <= 64'd36028797010575360;
            ROM0_arr[0][13] <= 64'd1;
            ROM0_arr[1][13] <= 64'd6366922389463153702;
            ROM0_arr[2][13] <= 64'd34359214072;
            ROM0_arr[3][13] <= 64'd8215369291935911999;
            ROM0_arr[4][13] <= 64'd18410715272404008961;
            ROM0_arr[5][13] <= 64'd17090085178304640863;
            ROM0_arr[6][13] <= 64'd288230376151710720;
            ROM0_arr[7][13] <= 64'd16192975500896648969;
            ROM0_arr[8][13] <= 64'd18446673700670423041;
            ROM0_arr[9][13] <= 64'd5834015391316509212;
            ROM0_arr[10][13] <= 64'd562949953421310;
            ROM0_arr[11][13] <= 64'd8930739766887302688;
            ROM0_arr[12][13] <= 64'd18446743931975630881;
            ROM0_arr[13][13] <= 64'd17449332314429639298;
            ROM0_arr[14][13] <= 64'd72058693532778496;
            ROM0_arr[15][13] <= 64'd17311265416183374564;
            ROM0_arr[0][14] <= 64'd1;
            ROM0_arr[1][14] <= 64'd288230376151712768;
            ROM0_arr[2][14] <= 64'd137438953440;
            ROM0_arr[3][14] <= 64'd140735340838912;
            ROM0_arr[4][14] <= 64'd18446739671368073217;
            ROM0_arr[5][14] <= 64'd18442240469787213841;
            ROM0_arr[6][14] <= 64'd32768;
            ROM0_arr[7][14] <= 64'd2199056809472;
            ROM0_arr[8][14] <= 64'd4503599626321920;
            ROM0_arr[9][14] <= 64'd4611615648609468416;
            ROM0_arr[10][14] <= 64'd18302628881338728449;
            ROM0_arr[11][14] <= 64'd18446744035055370249;
            ROM0_arr[12][14] <= 64'd1073741824;
            ROM0_arr[13][14] <= 64'd72058693532778496;
            ROM0_arr[14][14] <= 64'd18446744069414584313;
            ROM0_arr[15][14] <= 64'd16140901060200882177;
            ROM0_arr[0][15] <= 64'd1;
            ROM0_arr[1][15] <= 64'd9516004302527281633;
            ROM0_arr[2][15] <= 64'd274882101184;
            ROM0_arr[3][15] <= 64'd3341893669734556710;
            ROM0_arr[4][15] <= 64'd2305843008676823040;
            ROM0_arr[5][15] <= 64'd1116342470860912836;
            ROM0_arr[6][15] <= 64'd18446744035054321673;
            ROM0_arr[7][15] <= 64'd13417321343344118652;
            ROM0_arr[8][15] <= 64'd18158513693329981441;
            ROM0_arr[9][15] <= 64'd9083829225849678056;
            ROM0_arr[10][15] <= 64'd4295032831;
            ROM0_arr[11][15] <= 64'd7546206866789277329;
            ROM0_arr[12][15] <= 64'd36028797010575360;
            ROM0_arr[13][15] <= 64'd17311265416183374564;
            ROM0_arr[14][15] <= 64'd16140901060200882177;
            ROM0_arr[15][15] <= 64'd1362567150328163374;

            // ROM1 init
            ROM1_arr[0][0] <= 64'd1;
            ROM1_arr[1][0] <= 64'd1;
            ROM1_arr[2][0] <= 64'd1;
            ROM1_arr[3][0] <= 64'd1;
            ROM1_arr[4][0] <= 64'd1;
            ROM1_arr[5][0] <= 64'd1;
            ROM1_arr[6][0] <= 64'd1;
            ROM1_arr[7][0] <= 64'd1;
            ROM1_arr[8][0] <= 64'd1;
            ROM1_arr[9][0] <= 64'd1;
            ROM1_arr[10][0] <= 64'd1;
            ROM1_arr[11][0] <= 64'd1;
            ROM1_arr[12][0] <= 64'd1;
            ROM1_arr[13][0] <= 64'd1;
            ROM1_arr[14][0] <= 64'd1;
            ROM1_arr[15][0] <= 64'd1;
            ROM1_arr[0][1] <= 64'd1;
            ROM1_arr[1][1] <= 64'd14006830186316163511;
            ROM1_arr[2][1] <= 64'd15052656207385017564;
            ROM1_arr[3][1] <= 64'd9202451367179449552;
            ROM1_arr[4][1] <= 64'd1913039459307282826;
            ROM1_arr[5][1] <= 64'd10881114917016671572;
            ROM1_arr[6][1] <= 64'd10460593365646500703;
            ROM1_arr[7][1] <= 64'd3658040589001357399;
            ROM1_arr[8][1] <= 64'd12573252732142656207;
            ROM1_arr[9][1] <= 64'd13537781928143541450;
            ROM1_arr[10][1] <= 64'd7725134980519083461;
            ROM1_arr[11][1] <= 64'd15038653555595503587;
            ROM1_arr[12][1] <= 64'd15919780095311700439;
            ROM1_arr[13][1] <= 64'd3260171394465825874;
            ROM1_arr[14][1] <= 64'd14565379884206802520;
            ROM1_arr[15][1] <= 64'd16214251152771544261;
            ROM1_arr[0][2] <= 64'd1;
            ROM1_arr[1][2] <= 64'd15052656207385017564;
            ROM1_arr[2][2] <= 64'd1913039459307282826;
            ROM1_arr[3][2] <= 64'd10460593365646500703;
            ROM1_arr[4][2] <= 64'd12573252732142656207;
            ROM1_arr[5][2] <= 64'd7725134980519083461;
            ROM1_arr[6][2] <= 64'd15919780095311700439;
            ROM1_arr[7][2] <= 64'd14565379884206802520;
            ROM1_arr[8][2] <= 64'd11147770252432840497;
            ROM1_arr[9][2] <= 64'd11577486448795369550;
            ROM1_arr[10][2] <= 64'd11731715020642418612;
            ROM1_arr[11][2] <= 64'd12004140365210146681;
            ROM1_arr[12][2] <= 64'd6396200096592884887;
            ROM1_arr[13][2] <= 64'd8049782023765701561;
            ROM1_arr[14][2] <= 64'd12527349963958696492;
            ROM1_arr[15][2] <= 64'd3956111051294801955;
            ROM1_arr[0][3] <= 64'd1;
            ROM1_arr[1][3] <= 64'd9202451367179449552;
            ROM1_arr[2][3] <= 64'd10460593365646500703;
            ROM1_arr[3][3] <= 64'd13537781928143541450;
            ROM1_arr[4][3] <= 64'd15919780095311700439;
            ROM1_arr[5][3] <= 64'd16214251152771544261;
            ROM1_arr[6][3] <= 64'd11577486448795369550;
            ROM1_arr[7][3] <= 64'd14094041474627469271;
            ROM1_arr[8][3] <= 64'd6396200096592884887;
            ROM1_arr[9][3] <= 64'd3949970899253118150;
            ROM1_arr[10][3] <= 64'd3956111051294801955;
            ROM1_arr[11][3] <= 64'd3289556826179305825;
            ROM1_arr[12][3] <= 64'd8900146263973118671;
            ROM1_arr[13][3] <= 64'd9495908308903004412;
            ROM1_arr[14][3] <= 64'd17885125740710459782;
            ROM1_arr[15][3] <= 64'd7539172197244716846;
            ROM1_arr[0][4] <= 64'd1;
            ROM1_arr[1][4] <= 64'd1913039459307282826;
            ROM1_arr[2][4] <= 64'd12573252732142656207;
            ROM1_arr[3][4] <= 64'd15919780095311700439;
            ROM1_arr[4][4] <= 64'd11147770252432840497;
            ROM1_arr[5][4] <= 64'd11731715020642418612;
            ROM1_arr[6][4] <= 64'd6396200096592884887;
            ROM1_arr[7][4] <= 64'd12527349963958696492;
            ROM1_arr[8][4] <= 64'd18446181119461163011;
            ROM1_arr[9][4] <= 64'd8900146263973118671;
            ROM1_arr[10][4] <= 64'd15122929597976639421;
            ROM1_arr[11][4] <= 64'd2225341748615664720;
            ROM1_arr[12][4] <= 64'd6562114217670983589;
            ROM1_arr[13][4] <= 64'd7847524879092096009;
            ROM1_arr[14][4] <= 64'd875634265288439343;
            ROM1_arr[15][4] <= 64'd13440262264613344657;
            ROM1_arr[0][5] <= 64'd1;
            ROM1_arr[1][5] <= 64'd10881114917016671572;
            ROM1_arr[2][5] <= 64'd7725134980519083461;
            ROM1_arr[3][5] <= 64'd16214251152771544261;
            ROM1_arr[4][5] <= 64'd11731715020642418612;
            ROM1_arr[5][5] <= 64'd15646332241525257836;
            ROM1_arr[6][5] <= 64'd3956111051294801955;
            ROM1_arr[7][5] <= 64'd13566340103724003359;
            ROM1_arr[8][5] <= 64'd15122929597976639421;
            ROM1_arr[9][5] <= 64'd7539172197244716846;
            ROM1_arr[10][5] <= 64'd14091609828646341284;
            ROM1_arr[11][5] <= 64'd12882625803841659841;
            ROM1_arr[12][5] <= 64'd13440262264613344657;
            ROM1_arr[13][5] <= 64'd11784050230675421138;
            ROM1_arr[14][5] <= 64'd17516019197232489140;
            ROM1_arr[15][5] <= 64'd9443965423685914908;
            ROM1_arr[0][6] <= 64'd1;
            ROM1_arr[1][6] <= 64'd10460593365646500703;
            ROM1_arr[2][6] <= 64'd15919780095311700439;
            ROM1_arr[3][6] <= 64'd11577486448795369550;
            ROM1_arr[4][6] <= 64'd6396200096592884887;
            ROM1_arr[5][6] <= 64'd3956111051294801955;
            ROM1_arr[6][6] <= 64'd8900146263973118671;
            ROM1_arr[7][6] <= 64'd17885125740710459782;
            ROM1_arr[8][6] <= 64'd6562114217670983589;
            ROM1_arr[9][6] <= 64'd1305216586892671150;
            ROM1_arr[10][6] <= 64'd13440262264613344657;
            ROM1_arr[11][6] <= 64'd16182636211847971145;
            ROM1_arr[12][6] <= 64'd15245928743009060991;
            ROM1_arr[13][6] <= 64'd14885515920950843192;
            ROM1_arr[14][6] <= 64'd11323355628887372424;
            ROM1_arr[15][6] <= 64'd15089610673364298943;
            ROM1_arr[0][7] <= 64'd1;
            ROM1_arr[1][7] <= 64'd3658040589001357399;
            ROM1_arr[2][7] <= 64'd14565379884206802520;
            ROM1_arr[3][7] <= 64'd14094041474627469271;
            ROM1_arr[4][7] <= 64'd12527349963958696492;
            ROM1_arr[5][7] <= 64'd13566340103724003359;
            ROM1_arr[6][7] <= 64'd17885125740710459782;
            ROM1_arr[7][7] <= 64'd4065293009581645722;
            ROM1_arr[8][7] <= 64'd875634265288439343;
            ROM1_arr[9][7] <= 64'd10062399975831801284;
            ROM1_arr[10][7] <= 64'd17516019197232489140;
            ROM1_arr[11][7] <= 64'd4075317633252260392;
            ROM1_arr[12][7] <= 64'd11323355628887372424;
            ROM1_arr[13][7] <= 64'd17075652081414098800;
            ROM1_arr[14][7] <= 64'd12883701938510673118;
            ROM1_arr[15][7] <= 64'd2765937803960126615;
            ROM1_arr[0][8] <= 64'd1;
            ROM1_arr[1][8] <= 64'd12573252732142656207;
            ROM1_arr[2][8] <= 64'd11147770252432840497;
            ROM1_arr[3][8] <= 64'd6396200096592884887;
            ROM1_arr[4][8] <= 64'd18446181119461163011;
            ROM1_arr[5][8] <= 64'd15122929597976639421;
            ROM1_arr[6][8] <= 64'd6562114217670983589;
            ROM1_arr[7][8] <= 64'd875634265288439343;
            ROM1_arr[8][8] <= 64'd18444492269600899073;
            ROM1_arr[9][8] <= 64'd15245928743009060991;
            ROM1_arr[10][8] <= 64'd10853271128879547664;
            ROM1_arr[11][8] <= 64'd7673168496654431239;
            ROM1_arr[12][8] <= 64'd18442240469787213809;
            ROM1_arr[13][8] <= 64'd13787254465881465880;
            ROM1_arr[14][8] <= 64'd9362914843564906265;
            ROM1_arr[15][8] <= 64'd5240855794895625891;
            ROM1_arr[0][9] <= 64'd1;
            ROM1_arr[1][9] <= 64'd13537781928143541450;
            ROM1_arr[2][9] <= 64'd11577486448795369550;
            ROM1_arr[3][9] <= 64'd3949970899253118150;
            ROM1_arr[4][9] <= 64'd8900146263973118671;
            ROM1_arr[5][9] <= 64'd7539172197244716846;
            ROM1_arr[6][9] <= 64'd1305216586892671150;
            ROM1_arr[7][9] <= 64'd10062399975831801284;
            ROM1_arr[8][9] <= 64'd15245928743009060991;
            ROM1_arr[9][9] <= 64'd10140282184156893190;
            ROM1_arr[10][9] <= 64'd15089610673364298943;
            ROM1_arr[11][9] <= 64'd16966461843610068739;
            ROM1_arr[12][9] <= 64'd6431860813144680379;
            ROM1_arr[13][9] <= 64'd5209242550377892046;
            ROM1_arr[14][9] <= 64'd12590402701497627403;
            ROM1_arr[15][9] <= 64'd5693075206302722637;
            ROM1_arr[0][10] <= 64'd1;
            ROM1_arr[1][10] <= 64'd7725134980519083461;
            ROM1_arr[2][10] <= 64'd11731715020642418612;
            ROM1_arr[3][10] <= 64'd3956111051294801955;
            ROM1_arr[4][10] <= 64'd15122929597976639421;
            ROM1_arr[5][10] <= 64'd14091609828646341284;
            ROM1_arr[6][10] <= 64'd13440262264613344657;
            ROM1_arr[7][10] <= 64'd17516019197232489140;
            ROM1_arr[8][10] <= 64'd10853271128879547664;
            ROM1_arr[9][10] <= 64'd15089610673364298943;
            ROM1_arr[10][10] <= 64'd9983907413951898936;
            ROM1_arr[11][10] <= 64'd18085882527567857916;
            ROM1_arr[12][10] <= 64'd5240855794895625891;
            ROM1_arr[13][10] <= 64'd14307438406331844917;
            ROM1_arr[14][10] <= 64'd14151741787267893880;
            ROM1_arr[15][10] <= 64'd6498267541963153898;
            ROM1_arr[0][11] <= 64'd1;
            ROM1_arr[1][11] <= 64'd15038653555595503587;
            ROM1_arr[2][11] <= 64'd12004140365210146681;
            ROM1_arr[3][11] <= 64'd3289556826179305825;
            ROM1_arr[4][11] <= 64'd2225341748615664720;
            ROM1_arr[5][11] <= 64'd12882625803841659841;
            ROM1_arr[6][11] <= 64'd16182636211847971145;
            ROM1_arr[7][11] <= 64'd4075317633252260392;
            ROM1_arr[8][11] <= 64'd7673168496654431239;
            ROM1_arr[9][11] <= 64'd16966461843610068739;
            ROM1_arr[10][11] <= 64'd18085882527567857916;
            ROM1_arr[11][11] <= 64'd191154344862419240;
            ROM1_arr[12][11] <= 64'd6692683090235989383;
            ROM1_arr[13][11] <= 64'd13752338179252473593;
            ROM1_arr[14][11] <= 64'd1322784422603461084;
            ROM1_arr[15][11] <= 64'd6352413690540808131;
            ROM1_arr[0][12] <= 64'd1;
            ROM1_arr[1][12] <= 64'd15919780095311700439;
            ROM1_arr[2][12] <= 64'd6396200096592884887;
            ROM1_arr[3][12] <= 64'd8900146263973118671;
            ROM1_arr[4][12] <= 64'd6562114217670983589;
            ROM1_arr[5][12] <= 64'd13440262264613344657;
            ROM1_arr[6][12] <= 64'd15245928743009060991;
            ROM1_arr[7][12] <= 64'd11323355628887372424;
            ROM1_arr[8][12] <= 64'd18442240469787213809;
            ROM1_arr[9][12] <= 64'd6431860813144680379;
            ROM1_arr[10][12] <= 64'd5240855794895625891;
            ROM1_arr[11][12] <= 64'd6692683090235989383;
            ROM1_arr[12][12] <= 64'd5965722551466996711;
            ROM1_arr[13][12] <= 64'd9906341360885134636;
            ROM1_arr[14][12] <= 64'd9809941408468046069;
            ROM1_arr[15][12] <= 64'd14267241681714216412;
            ROM1_arr[0][13] <= 64'd1;
            ROM1_arr[1][13] <= 64'd3260171394465825874;
            ROM1_arr[2][13] <= 64'd8049782023765701561;
            ROM1_arr[3][13] <= 64'd9495908308903004412;
            ROM1_arr[4][13] <= 64'd7847524879092096009;
            ROM1_arr[5][13] <= 64'd11784050230675421138;
            ROM1_arr[6][13] <= 64'd14885515920950843192;
            ROM1_arr[7][13] <= 64'd17075652081414098800;
            ROM1_arr[8][13] <= 64'd13787254465881465880;
            ROM1_arr[9][13] <= 64'd5209242550377892046;
            ROM1_arr[10][13] <= 64'd14307438406331844917;
            ROM1_arr[11][13] <= 64'd13752338179252473593;
            ROM1_arr[12][13] <= 64'd9906341360885134636;
            ROM1_arr[13][13] <= 64'd17081697152343396870;
            ROM1_arr[14][13] <= 64'd8699858785941968005;
            ROM1_arr[15][13] <= 64'd2740180791756161213;
            ROM1_arr[0][14] <= 64'd1;
            ROM1_arr[1][14] <= 64'd14565379884206802520;
            ROM1_arr[2][14] <= 64'd12527349963958696492;
            ROM1_arr[3][14] <= 64'd17885125740710459782;
            ROM1_arr[4][14] <= 64'd875634265288439343;
            ROM1_arr[5][14] <= 64'd17516019197232489140;
            ROM1_arr[6][14] <= 64'd11323355628887372424;
            ROM1_arr[7][14] <= 64'd12883701938510673118;
            ROM1_arr[8][14] <= 64'd9362914843564906265;
            ROM1_arr[9][14] <= 64'd12590402701497627403;
            ROM1_arr[10][14] <= 64'd14151741787267893880;
            ROM1_arr[11][14] <= 64'd1322784422603461084;
            ROM1_arr[12][14] <= 64'd9809941408468046069;
            ROM1_arr[13][14] <= 64'd8699858785941968005;
            ROM1_arr[14][14] <= 64'd10757588516645913927;
            ROM1_arr[15][14] <= 64'd14377936972942800771;
            ROM1_arr[0][15] <= 64'd1;
            ROM1_arr[1][15] <= 64'd16214251152771544261;
            ROM1_arr[2][15] <= 64'd3956111051294801955;
            ROM1_arr[3][15] <= 64'd7539172197244716846;
            ROM1_arr[4][15] <= 64'd13440262264613344657;
            ROM1_arr[5][15] <= 64'd9443965423685914908;
            ROM1_arr[6][15] <= 64'd15089610673364298943;
            ROM1_arr[7][15] <= 64'd2765937803960126615;
            ROM1_arr[8][15] <= 64'd5240855794895625891;
            ROM1_arr[9][15] <= 64'd5693075206302722637;
            ROM1_arr[10][15] <= 64'd6498267541963153898;
            ROM1_arr[11][15] <= 64'd6352413690540808131;
            ROM1_arr[12][15] <= 64'd14267241681714216412;
            ROM1_arr[13][15] <= 64'd2740180791756161213;
            ROM1_arr[14][15] <= 64'd14377936972942800771;
            ROM1_arr[15][15] <= 64'd14148553018161426505;
            // ROM2 init
            ROM2_arr[0][0] <= 64'd1;
            ROM2_arr[1][0] <= 64'd1;
            ROM2_arr[2][0] <= 64'd1;
            ROM2_arr[3][0] <= 64'd1;
            ROM2_arr[4][0] <= 64'd1;
            ROM2_arr[5][0] <= 64'd1;
            ROM2_arr[6][0] <= 64'd1;
            ROM2_arr[7][0] <= 64'd1;
            ROM2_arr[8][0] <= 64'd1;
            ROM2_arr[9][0] <= 64'd1;
            ROM2_arr[10][0] <= 64'd1;
            ROM2_arr[11][0] <= 64'd1;
            ROM2_arr[12][0] <= 64'd1;
            ROM2_arr[13][0] <= 64'd1;
            ROM2_arr[14][0] <= 64'd1;
            ROM2_arr[15][0] <= 64'd1;
            ROM2_arr[0][1] <= 64'd1;
            ROM2_arr[1][1] <= 64'd14603442835287214144;
            ROM2_arr[2][1] <= 64'd14092008124193502130;
            ROM2_arr[3][1] <= 64'd6886462153987203820;
            ROM2_arr[4][1] <= 64'd4043556811946972802;
            ROM2_arr[5][1] <= 64'd2840400505270878937;
            ROM2_arr[6][1] <= 64'd18138845337817616439;
            ROM2_arr[7][1] <= 64'd9927864368106092497;
            ROM2_arr[8][1] <= 64'd9071165522957276205;
            ROM2_arr[9][1] <= 64'd2655872976626746565;
            ROM2_arr[10][1] <= 64'd11703777381874358041;
            ROM2_arr[11][1] <= 64'd7492191627268029833;
            ROM2_arr[12][1] <= 64'd10474213472750683764;
            ROM2_arr[13][1] <= 64'd5020150431739777697;
            ROM2_arr[14][1] <= 64'd16666718547735378570;
            ROM2_arr[15][1] <= 64'd16433623054813571938;
            ROM2_arr[0][2] <= 64'd1;
            ROM2_arr[1][2] <= 64'd14092008124193502130;
            ROM2_arr[2][2] <= 64'd4043556811946972802;
            ROM2_arr[3][2] <= 64'd18138845337817616439;
            ROM2_arr[4][2] <= 64'd9071165522957276205;
            ROM2_arr[5][2] <= 64'd11703777381874358041;
            ROM2_arr[6][2] <= 64'd10474213472750683764;
            ROM2_arr[7][2] <= 64'd16666718547735378570;
            ROM2_arr[8][2] <= 64'd14006830186316163511;
            ROM2_arr[9][2] <= 64'd18414194918738960790;
            ROM2_arr[10][2] <= 64'd2676548733418181014;
            ROM2_arr[11][2] <= 64'd17231931100285778307;
            ROM2_arr[12][2] <= 64'd2452125344670730664;
            ROM2_arr[13][2] <= 64'd17561784851306960425;
            ROM2_arr[14][2] <= 64'd15529017648405328904;
            ROM2_arr[15][2] <= 64'd11433841022347624621;
            ROM2_arr[0][3] <= 64'd1;
            ROM2_arr[1][3] <= 64'd6886462153987203820;
            ROM2_arr[2][3] <= 64'd18138845337817616439;
            ROM2_arr[3][3] <= 64'd2655872976626746565;
            ROM2_arr[4][3] <= 64'd10474213472750683764;
            ROM2_arr[5][3] <= 64'd16433623054813571938;
            ROM2_arr[6][3] <= 64'd18414194918738960790;
            ROM2_arr[7][3] <= 64'd12089335110147162665;
            ROM2_arr[8][3] <= 64'd2452125344670730664;
            ROM2_arr[9][3] <= 64'd14620677213708548715;
            ROM2_arr[10][3] <= 64'd11433841022347624621;
            ROM2_arr[11][3] <= 64'd6269618961335635998;
            ROM2_arr[12][3] <= 64'd5350167283985131626;
            ROM2_arr[13][3] <= 64'd11077481226347603699;
            ROM2_arr[14][3] <= 64'd3792960320742134233;
            ROM2_arr[15][3] <= 64'd6767729679576688768;
            ROM2_arr[0][4] <= 64'd1;
            ROM2_arr[1][4] <= 64'd4043556811946972802;
            ROM2_arr[2][4] <= 64'd9071165522957276205;
            ROM2_arr[3][4] <= 64'd10474213472750683764;
            ROM2_arr[4][4] <= 64'd14006830186316163511;
            ROM2_arr[5][4] <= 64'd2676548733418181014;
            ROM2_arr[6][4] <= 64'd2452125344670730664;
            ROM2_arr[7][4] <= 64'd15529017648405328904;
            ROM2_arr[8][4] <= 64'd15052656207385017564;
            ROM2_arr[9][4] <= 64'd5350167283985131626;
            ROM2_arr[10][4] <= 64'd638849890512999907;
            ROM2_arr[11][4] <= 64'd3292571118866816134;
            ROM2_arr[12][4] <= 64'd9202451367179449552;
            ROM2_arr[13][4] <= 64'd8487349938101489318;
            ROM2_arr[14][4] <= 64'd537896514274431823;
            ROM2_arr[15][4] <= 64'd7734123025605687877;
            ROM2_arr[0][5] <= 64'd1;
            ROM2_arr[1][5] <= 64'd2840400505270878937;
            ROM2_arr[2][5] <= 64'd11703777381874358041;
            ROM2_arr[3][5] <= 64'd16433623054813571938;
            ROM2_arr[4][5] <= 64'd2676548733418181014;
            ROM2_arr[5][5] <= 64'd8858629302739700209;
            ROM2_arr[6][5] <= 64'd11433841022347624621;
            ROM2_arr[7][5] <= 64'd10148874914461315166;
            ROM2_arr[8][5] <= 64'd638849890512999907;
            ROM2_arr[9][5] <= 64'd6767729679576688768;
            ROM2_arr[10][5] <= 64'd16462828118252960335;
            ROM2_arr[11][5] <= 64'd16721623190635630841;
            ROM2_arr[12][5] <= 64'd7734123025605687877;
            ROM2_arr[13][5] <= 64'd14702451440905515216;
            ROM2_arr[14][5] <= 64'd2775966812770153583;
            ROM2_arr[15][5] <= 64'd16803758761047781263;
            ROM2_arr[0][6] <= 64'd1;
            ROM2_arr[1][6] <= 64'd18138845337817616439;
            ROM2_arr[2][6] <= 64'd10474213472750683764;
            ROM2_arr[3][6] <= 64'd18414194918738960790;
            ROM2_arr[4][6] <= 64'd2452125344670730664;
            ROM2_arr[5][6] <= 64'd11433841022347624621;
            ROM2_arr[6][6] <= 64'd5350167283985131626;
            ROM2_arr[7][6] <= 64'd3792960320742134233;
            ROM2_arr[8][6] <= 64'd9202451367179449552;
            ROM2_arr[9][6] <= 64'd12450734428395028578;
            ROM2_arr[10][6] <= 64'd7734123025605687877;
            ROM2_arr[11][6] <= 64'd17491778934546556896;
            ROM2_arr[12][6] <= 64'd15583913849859751243;
            ROM2_arr[13][6] <= 64'd11527892611242128361;
            ROM2_arr[14][6] <= 64'd283879498861853653;
            ROM2_arr[15][6] <= 64'd418570971427346365;
            ROM2_arr[0][7] <= 64'd1;
            ROM2_arr[1][7] <= 64'd9927864368106092497;
            ROM2_arr[2][7] <= 64'd16666718547735378570;
            ROM2_arr[3][7] <= 64'd12089335110147162665;
            ROM2_arr[4][7] <= 64'd15529017648405328904;
            ROM2_arr[5][7] <= 64'd10148874914461315166;
            ROM2_arr[6][7] <= 64'd3792960320742134233;
            ROM2_arr[7][7] <= 64'd624304266358974706;
            ROM2_arr[8][7] <= 64'd537896514274431823;
            ROM2_arr[9][7] <= 64'd4049320560851992053;
            ROM2_arr[10][7] <= 64'd2775966812770153583;
            ROM2_arr[11][7] <= 64'd601746077641686379;
            ROM2_arr[12][7] <= 64'd283879498861853653;
            ROM2_arr[13][7] <= 64'd15937576857968480300;
            ROM2_arr[14][7] <= 64'd9854506929839881396;
            ROM2_arr[15][7] <= 64'd14654049273797424740;
            ROM2_arr[0][8] <= 64'd1;
            ROM2_arr[1][8] <= 64'd9071165522957276205;
            ROM2_arr[2][8] <= 64'd14006830186316163511;
            ROM2_arr[3][8] <= 64'd2452125344670730664;
            ROM2_arr[4][8] <= 64'd15052656207385017564;
            ROM2_arr[5][8] <= 64'd638849890512999907;
            ROM2_arr[6][8] <= 64'd9202451367179449552;
            ROM2_arr[7][8] <= 64'd537896514274431823;
            ROM2_arr[8][8] <= 64'd1913039459307282826;
            ROM2_arr[9][8] <= 64'd15583913849859751243;
            ROM2_arr[10][8] <= 64'd10881114917016671572;
            ROM2_arr[11][8] <= 64'd172919261666014791;
            ROM2_arr[12][8] <= 64'd10460593365646500703;
            ROM2_arr[13][8] <= 64'd17572224462131996077;
            ROM2_arr[14][8] <= 64'd3658040589001357399;
            ROM2_arr[15][8] <= 64'd11260516089836515982;
            ROM2_arr[0][9] <= 64'd1;
            ROM2_arr[1][9] <= 64'd2655872976626746565;
            ROM2_arr[2][9] <= 64'd18414194918738960790;
            ROM2_arr[3][9] <= 64'd14620677213708548715;
            ROM2_arr[4][9] <= 64'd5350167283985131626;
            ROM2_arr[5][9] <= 64'd6767729679576688768;
            ROM2_arr[6][9] <= 64'd12450734428395028578;
            ROM2_arr[7][9] <= 64'd4049320560851992053;
            ROM2_arr[8][9] <= 64'd15583913849859751243;
            ROM2_arr[9][9] <= 64'd7758667811057267014;
            ROM2_arr[10][9] <= 64'd418570971427346365;
            ROM2_arr[11][9] <= 64'd16096405968772420831;
            ROM2_arr[12][9] <= 64'd17577632102214582396;
            ROM2_arr[13][9] <= 64'd18120918623894693431;
            ROM2_arr[14][9] <= 64'd12344405285182455956;
            ROM2_arr[15][9] <= 64'd974417746440743327;
            ROM2_arr[0][10] <= 64'd1;
            ROM2_arr[1][10] <= 64'd11703777381874358041;
            ROM2_arr[2][10] <= 64'd2676548733418181014;
            ROM2_arr[3][10] <= 64'd11433841022347624621;
            ROM2_arr[4][10] <= 64'd638849890512999907;
            ROM2_arr[5][10] <= 64'd16462828118252960335;
            ROM2_arr[6][10] <= 64'd7734123025605687877;
            ROM2_arr[7][10] <= 64'd2775966812770153583;
            ROM2_arr[8][10] <= 64'd10881114917016671572;
            ROM2_arr[9][10] <= 64'd418570971427346365;
            ROM2_arr[10][10] <= 64'd11888488389018040474;
            ROM2_arr[11][10] <= 64'd10881384902014718835;
            ROM2_arr[12][10] <= 64'd11260516089836515982;
            ROM2_arr[13][10] <= 64'd5511237480569377606;
            ROM2_arr[14][10] <= 64'd13253372258298764714;
            ROM2_arr[15][10] <= 64'd2443842004063759267;
            ROM2_arr[0][11] <= 64'd1;
            ROM2_arr[1][11] <= 64'd7492191627268029833;
            ROM2_arr[2][11] <= 64'd17231931100285778307;
            ROM2_arr[3][11] <= 64'd6269618961335635998;
            ROM2_arr[4][11] <= 64'd3292571118866816134;
            ROM2_arr[5][11] <= 64'd16721623190635630841;
            ROM2_arr[6][11] <= 64'd17491778934546556896;
            ROM2_arr[7][11] <= 64'd601746077641686379;
            ROM2_arr[8][11] <= 64'd172919261666014791;
            ROM2_arr[9][11] <= 64'd16096405968772420831;
            ROM2_arr[10][11] <= 64'd10881384902014718835;
            ROM2_arr[11][11] <= 64'd12222620110109638483;
            ROM2_arr[12][11] <= 64'd15395467146316174056;
            ROM2_arr[13][11] <= 64'd7403481904734983592;
            ROM2_arr[14][11] <= 64'd9667434717573275621;
            ROM2_arr[15][11] <= 64'd9314406845994532780;
            ROM2_arr[0][12] <= 64'd1;
            ROM2_arr[1][12] <= 64'd10474213472750683764;
            ROM2_arr[2][12] <= 64'd2452125344670730664;
            ROM2_arr[3][12] <= 64'd5350167283985131626;
            ROM2_arr[4][12] <= 64'd9202451367179449552;
            ROM2_arr[5][12] <= 64'd7734123025605687877;
            ROM2_arr[6][12] <= 64'd15583913849859751243;
            ROM2_arr[7][12] <= 64'd283879498861853653;
            ROM2_arr[8][12] <= 64'd10460593365646500703;
            ROM2_arr[9][12] <= 64'd17577632102214582396;
            ROM2_arr[10][12] <= 64'd11260516089836515982;
            ROM2_arr[11][12] <= 64'd15395467146316174056;
            ROM2_arr[12][12] <= 64'd13537781928143541450;
            ROM2_arr[13][12] <= 64'd6295673273103589313;
            ROM2_arr[14][12] <= 64'd13606998934696871123;
            ROM2_arr[15][12] <= 64'd13069618832511821766;
            ROM2_arr[0][13] <= 64'd1;
            ROM2_arr[1][13] <= 64'd5020150431739777697;
            ROM2_arr[2][13] <= 64'd17561784851306960425;
            ROM2_arr[3][13] <= 64'd11077481226347603699;
            ROM2_arr[4][13] <= 64'd8487349938101489318;
            ROM2_arr[5][13] <= 64'd14702451440905515216;
            ROM2_arr[6][13] <= 64'd11527892611242128361;
            ROM2_arr[7][13] <= 64'd15937576857968480300;
            ROM2_arr[8][13] <= 64'd17572224462131996077;
            ROM2_arr[9][13] <= 64'd18120918623894693431;
            ROM2_arr[10][13] <= 64'd5511237480569377606;
            ROM2_arr[11][13] <= 64'd7403481904734983592;
            ROM2_arr[12][13] <= 64'd6295673273103589313;
            ROM2_arr[13][13] <= 64'd4058470387566679753;
            ROM2_arr[14][13] <= 64'd803938878720571184;
            ROM2_arr[15][13] <= 64'd11695028341473597159;
            ROM2_arr[0][14] <= 64'd1;
            ROM2_arr[1][14] <= 64'd16666718547735378570;
            ROM2_arr[2][14] <= 64'd15529017648405328904;
            ROM2_arr[3][14] <= 64'd3792960320742134233;
            ROM2_arr[4][14] <= 64'd537896514274431823;
            ROM2_arr[5][14] <= 64'd2775966812770153583;
            ROM2_arr[6][14] <= 64'd283879498861853653;
            ROM2_arr[7][14] <= 64'd9854506929839881396;
            ROM2_arr[8][14] <= 64'd3658040589001357399;
            ROM2_arr[9][14] <= 64'd12344405285182455956;
            ROM2_arr[10][14] <= 64'd13253372258298764714;
            ROM2_arr[11][14] <= 64'd9667434717573275621;
            ROM2_arr[12][14] <= 64'd13606998934696871123;
            ROM2_arr[13][14] <= 64'd803938878720571184;
            ROM2_arr[14][14] <= 64'd12358063764579062105;
            ROM2_arr[15][14] <= 64'd16630061566374667835;
            ROM2_arr[0][15] <= 64'd1;
            ROM2_arr[1][15] <= 64'd16433623054813571938;
            ROM2_arr[2][15] <= 64'd11433841022347624621;
            ROM2_arr[3][15] <= 64'd6767729679576688768;
            ROM2_arr[4][15] <= 64'd7734123025605687877;
            ROM2_arr[5][15] <= 64'd16803758761047781263;
            ROM2_arr[6][15] <= 64'd418570971427346365;
            ROM2_arr[7][15] <= 64'd14654049273797424740;
            ROM2_arr[8][15] <= 64'd11260516089836515982;
            ROM2_arr[9][15] <= 64'd974417746440743327;
            ROM2_arr[10][15] <= 64'd2443842004063759267;
            ROM2_arr[11][15] <= 64'd9314406845994532780;
            ROM2_arr[12][15] <= 64'd13069618832511821766;
            ROM2_arr[13][15] <= 64'd11695028341473597159;
            ROM2_arr[14][15] <= 64'd16630061566374667835;
            ROM2_arr[15][15] <= 64'd9158626267514805997;
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM0_b0     <= 64'd0    ;
            ROM0_b1     <= 64'd0    ;
            ROM0_b2     <= 64'd0    ;
            ROM0_b3     <= 64'd0    ;
            ROM0_b4     <= 64'd0    ;
            ROM0_b5     <= 64'd0    ;
            ROM0_b6     <= 64'd0    ;
            ROM0_b7     <= 64'd0    ;
            ROM0_b8     <= 64'd0    ;
            ROM0_b9     <= 64'd0    ;
            ROM0_b10    <= 64'd0    ;
            ROM0_b11    <= 64'd0    ;
            ROM0_b12    <= 64'd0    ; 
            ROM0_b13    <= 64'd0    ;
            ROM0_b14    <= 64'd0    ; 
            ROM0_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (MA0)
                    4'd0:
                        begin
                            ROM0_b0     <=  ROM0_arr[0][0]  ;
                            ROM0_b1     <=  ROM0_arr[0][1]  ;
                            ROM0_b2     <=  ROM0_arr[0][2]  ;
                            ROM0_b3     <=  ROM0_arr[0][3]  ;
                            ROM0_b4     <=  ROM0_arr[0][4]  ;
                            ROM0_b5     <=  ROM0_arr[0][5]  ;
                            ROM0_b6     <=  ROM0_arr[0][6]  ;
                            ROM0_b7     <=  ROM0_arr[0][7]  ;
                            ROM0_b8     <=  ROM0_arr[0][8]  ;
                            ROM0_b9     <=  ROM0_arr[0][9]  ;
                            ROM0_b10    <=  ROM0_arr[0][10] ;
                            ROM0_b11    <=  ROM0_arr[0][11] ;
                            ROM0_b12    <=  ROM0_arr[0][12] ;
                            ROM0_b13    <=  ROM0_arr[0][13] ;
                            ROM0_b14    <=  ROM0_arr[0][14] ;
                            ROM0_b15    <=  ROM0_arr[0][15] ;
                        end
                    4'd1:
                        begin
                            ROM0_b0     <=  ROM0_arr[1][0]  ;
                            ROM0_b1     <=  ROM0_arr[1][1]  ;
                            ROM0_b2     <=  ROM0_arr[1][2]  ;
                            ROM0_b3     <=  ROM0_arr[1][3]  ;
                            ROM0_b4     <=  ROM0_arr[1][4]  ;
                            ROM0_b5     <=  ROM0_arr[1][5]  ;
                            ROM0_b6     <=  ROM0_arr[1][6]  ;
                            ROM0_b7     <=  ROM0_arr[1][7]  ;
                            ROM0_b8     <=  ROM0_arr[1][8]  ;
                            ROM0_b9     <=  ROM0_arr[1][9]  ;
                            ROM0_b10    <=  ROM0_arr[1][10] ;
                            ROM0_b11    <=  ROM0_arr[1][11] ;
                            ROM0_b12    <=  ROM0_arr[1][12] ;
                            ROM0_b13    <=  ROM0_arr[1][13] ;
                            ROM0_b14    <=  ROM0_arr[1][14] ;
                            ROM0_b15    <=  ROM0_arr[1][15] ;
                        end
                    4'd2:
                        begin
                            ROM0_b0     <=  ROM0_arr[2][0]  ;
                            ROM0_b1     <=  ROM0_arr[2][1]  ;
                            ROM0_b2     <=  ROM0_arr[2][2]  ;
                            ROM0_b3     <=  ROM0_arr[2][3]  ;
                            ROM0_b4     <=  ROM0_arr[2][4]  ;
                            ROM0_b5     <=  ROM0_arr[2][5]  ;
                            ROM0_b6     <=  ROM0_arr[2][6]  ;
                            ROM0_b7     <=  ROM0_arr[2][7]  ;
                            ROM0_b8     <=  ROM0_arr[2][8]  ;
                            ROM0_b9     <=  ROM0_arr[2][9]  ;
                            ROM0_b10    <=  ROM0_arr[2][10] ;
                            ROM0_b11    <=  ROM0_arr[2][11] ;
                            ROM0_b12    <=  ROM0_arr[2][12] ;
                            ROM0_b13    <=  ROM0_arr[2][13] ;
                            ROM0_b14    <=  ROM0_arr[2][14] ;
                            ROM0_b15    <=  ROM0_arr[2][15] ;
                        end
                    4'd3:
                        begin
                            ROM0_b0     <=  ROM0_arr[3][0]  ;
                            ROM0_b1     <=  ROM0_arr[3][1]  ;
                            ROM0_b2     <=  ROM0_arr[3][2]  ;
                            ROM0_b3     <=  ROM0_arr[3][3]  ;
                            ROM0_b4     <=  ROM0_arr[3][4]  ;
                            ROM0_b5     <=  ROM0_arr[3][5]  ;
                            ROM0_b6     <=  ROM0_arr[3][6]  ;
                            ROM0_b7     <=  ROM0_arr[3][7]  ;
                            ROM0_b8     <=  ROM0_arr[3][8]  ;
                            ROM0_b9     <=  ROM0_arr[3][9]  ;
                            ROM0_b10    <=  ROM0_arr[3][10] ;
                            ROM0_b11    <=  ROM0_arr[3][11] ;
                            ROM0_b12    <=  ROM0_arr[3][12] ;
                            ROM0_b13    <=  ROM0_arr[3][13] ;
                            ROM0_b14    <=  ROM0_arr[3][14] ;
                            ROM0_b15    <=  ROM0_arr[3][15] ;
                        end
                    4'd4:
                        begin
                            ROM0_b0     <=  ROM0_arr[4][0]  ;
                            ROM0_b1     <=  ROM0_arr[4][1]  ;
                            ROM0_b2     <=  ROM0_arr[4][2]  ;
                            ROM0_b3     <=  ROM0_arr[4][3]  ;
                            ROM0_b4     <=  ROM0_arr[4][4]  ;
                            ROM0_b5     <=  ROM0_arr[4][5]  ;
                            ROM0_b6     <=  ROM0_arr[4][6]  ;
                            ROM0_b7     <=  ROM0_arr[4][7]  ;
                            ROM0_b8     <=  ROM0_arr[4][8]  ;
                            ROM0_b9     <=  ROM0_arr[4][9]  ;
                            ROM0_b10    <=  ROM0_arr[4][10] ;
                            ROM0_b11    <=  ROM0_arr[4][11] ;
                            ROM0_b12    <=  ROM0_arr[4][12] ;
                            ROM0_b13    <=  ROM0_arr[4][13] ;
                            ROM0_b14    <=  ROM0_arr[4][14] ;
                            ROM0_b15    <=  ROM0_arr[4][15] ;
                        end
                    4'd5:
                        begin
                            ROM0_b0     <=  ROM0_arr[5][0]  ;
                            ROM0_b1     <=  ROM0_arr[5][1]  ;
                            ROM0_b2     <=  ROM0_arr[5][2]  ;
                            ROM0_b3     <=  ROM0_arr[5][3]  ;
                            ROM0_b4     <=  ROM0_arr[5][4]  ;
                            ROM0_b5     <=  ROM0_arr[5][5]  ;
                            ROM0_b6     <=  ROM0_arr[5][6]  ;
                            ROM0_b7     <=  ROM0_arr[5][7]  ;
                            ROM0_b8     <=  ROM0_arr[5][8]  ;
                            ROM0_b9     <=  ROM0_arr[5][9]  ;
                            ROM0_b10    <=  ROM0_arr[5][10] ;
                            ROM0_b11    <=  ROM0_arr[5][11] ;
                            ROM0_b12    <=  ROM0_arr[5][12] ;
                            ROM0_b13    <=  ROM0_arr[5][13] ;
                            ROM0_b14    <=  ROM0_arr[5][14] ;
                            ROM0_b15    <=  ROM0_arr[5][15] ;
                        end
                    4'd6:
                        begin
                            ROM0_b0     <=  ROM0_arr[6][0]  ;
                            ROM0_b1     <=  ROM0_arr[6][1]  ;
                            ROM0_b2     <=  ROM0_arr[6][2]  ;
                            ROM0_b3     <=  ROM0_arr[6][3]  ;
                            ROM0_b4     <=  ROM0_arr[6][4]  ;
                            ROM0_b5     <=  ROM0_arr[6][5]  ;
                            ROM0_b6     <=  ROM0_arr[6][6]  ;
                            ROM0_b7     <=  ROM0_arr[6][7]  ;
                            ROM0_b8     <=  ROM0_arr[6][8]  ;
                            ROM0_b9     <=  ROM0_arr[6][9]  ;
                            ROM0_b10    <=  ROM0_arr[6][10] ;
                            ROM0_b11    <=  ROM0_arr[6][11] ;
                            ROM0_b12    <=  ROM0_arr[6][12] ;
                            ROM0_b13    <=  ROM0_arr[6][13] ;
                            ROM0_b14    <=  ROM0_arr[6][14] ;
                            ROM0_b15    <=  ROM0_arr[6][15] ;
                        end
                    4'd7:
                        begin
                            ROM0_b0     <=  ROM0_arr[7][0]  ;
                            ROM0_b1     <=  ROM0_arr[7][1]  ;
                            ROM0_b2     <=  ROM0_arr[7][2]  ;
                            ROM0_b3     <=  ROM0_arr[7][3]  ;
                            ROM0_b4     <=  ROM0_arr[7][4]  ;
                            ROM0_b5     <=  ROM0_arr[7][5]  ;
                            ROM0_b6     <=  ROM0_arr[7][6]  ;
                            ROM0_b7     <=  ROM0_arr[7][7]  ;
                            ROM0_b8     <=  ROM0_arr[7][8]  ;
                            ROM0_b9     <=  ROM0_arr[7][9]  ;
                            ROM0_b10    <=  ROM0_arr[7][10] ;
                            ROM0_b11    <=  ROM0_arr[7][11] ;
                            ROM0_b12    <=  ROM0_arr[7][12] ;
                            ROM0_b13    <=  ROM0_arr[7][13] ;
                            ROM0_b14    <=  ROM0_arr[7][14] ;
                            ROM0_b15    <=  ROM0_arr[7][15] ;
                        end
                    4'd8:
                        begin
                            ROM0_b0     <=  ROM0_arr[8][0]  ;
                            ROM0_b1     <=  ROM0_arr[8][1]  ;
                            ROM0_b2     <=  ROM0_arr[8][2]  ;
                            ROM0_b3     <=  ROM0_arr[8][3]  ;
                            ROM0_b4     <=  ROM0_arr[8][4]  ;
                            ROM0_b5     <=  ROM0_arr[8][5]  ;
                            ROM0_b6     <=  ROM0_arr[8][6]  ;
                            ROM0_b7     <=  ROM0_arr[8][7]  ;
                            ROM0_b8     <=  ROM0_arr[8][8]  ;
                            ROM0_b9     <=  ROM0_arr[8][9]  ;
                            ROM0_b10    <=  ROM0_arr[8][10] ;
                            ROM0_b11    <=  ROM0_arr[8][11] ;
                            ROM0_b12    <=  ROM0_arr[8][12] ;
                            ROM0_b13    <=  ROM0_arr[8][13] ;
                            ROM0_b14    <=  ROM0_arr[8][14] ;
                            ROM0_b15    <=  ROM0_arr[8][15] ;
                        end
                    4'd9:
                        begin
                            ROM0_b0     <=  ROM0_arr[9][0]  ;
                            ROM0_b1     <=  ROM0_arr[9][1]  ;
                            ROM0_b2     <=  ROM0_arr[9][2]  ;
                            ROM0_b3     <=  ROM0_arr[9][3]  ;
                            ROM0_b4     <=  ROM0_arr[9][4]  ;
                            ROM0_b5     <=  ROM0_arr[9][5]  ;
                            ROM0_b6     <=  ROM0_arr[9][6]  ;
                            ROM0_b7     <=  ROM0_arr[9][7]  ;
                            ROM0_b8     <=  ROM0_arr[9][8]  ;
                            ROM0_b9     <=  ROM0_arr[9][9]  ;
                            ROM0_b10    <=  ROM0_arr[9][10] ;
                            ROM0_b11    <=  ROM0_arr[9][11] ;
                            ROM0_b12    <=  ROM0_arr[9][12] ;
                            ROM0_b13    <=  ROM0_arr[9][13] ;
                            ROM0_b14    <=  ROM0_arr[9][14] ;
                            ROM0_b15    <=  ROM0_arr[9][15] ;
                        end
                    4'd10:
                        begin
                            ROM0_b0     <=  ROM0_arr[10][0]  ;
                            ROM0_b1     <=  ROM0_arr[10][1]  ;
                            ROM0_b2     <=  ROM0_arr[10][2]  ;
                            ROM0_b3     <=  ROM0_arr[10][3]  ;
                            ROM0_b4     <=  ROM0_arr[10][4]  ;
                            ROM0_b5     <=  ROM0_arr[10][5]  ;
                            ROM0_b6     <=  ROM0_arr[10][6]  ;
                            ROM0_b7     <=  ROM0_arr[10][7]  ;
                            ROM0_b8     <=  ROM0_arr[10][8]  ;
                            ROM0_b9     <=  ROM0_arr[10][9]  ;
                            ROM0_b10    <=  ROM0_arr[10][10] ;
                            ROM0_b11    <=  ROM0_arr[10][11] ;
                            ROM0_b12    <=  ROM0_arr[10][12] ;
                            ROM0_b13    <=  ROM0_arr[10][13] ;
                            ROM0_b14    <=  ROM0_arr[10][14] ;
                            ROM0_b15    <=  ROM0_arr[10][15] ;
                        end
                    4'd11:
                        begin
                            ROM0_b0     <=  ROM0_arr[11][0]  ;
                            ROM0_b1     <=  ROM0_arr[11][1]  ;
                            ROM0_b2     <=  ROM0_arr[11][2]  ;
                            ROM0_b3     <=  ROM0_arr[11][3]  ;
                            ROM0_b4     <=  ROM0_arr[11][4]  ;
                            ROM0_b5     <=  ROM0_arr[11][5]  ;
                            ROM0_b6     <=  ROM0_arr[11][6]  ;
                            ROM0_b7     <=  ROM0_arr[11][7]  ;
                            ROM0_b8     <=  ROM0_arr[11][8]  ;
                            ROM0_b9     <=  ROM0_arr[11][9]  ;
                            ROM0_b10    <=  ROM0_arr[11][10] ;
                            ROM0_b11    <=  ROM0_arr[11][11] ;
                            ROM0_b12    <=  ROM0_arr[11][12] ;
                            ROM0_b13    <=  ROM0_arr[11][13] ;
                            ROM0_b14    <=  ROM0_arr[11][14] ;
                            ROM0_b15    <=  ROM0_arr[11][15] ;
                        end
                    4'd12:
                        begin
                            ROM0_b0     <=  ROM0_arr[12][0]  ;
                            ROM0_b1     <=  ROM0_arr[12][1]  ;
                            ROM0_b2     <=  ROM0_arr[12][2]  ;
                            ROM0_b3     <=  ROM0_arr[12][3]  ;
                            ROM0_b4     <=  ROM0_arr[12][4]  ;
                            ROM0_b5     <=  ROM0_arr[12][5]  ;
                            ROM0_b6     <=  ROM0_arr[12][6]  ;
                            ROM0_b7     <=  ROM0_arr[12][7]  ;
                            ROM0_b8     <=  ROM0_arr[12][8]  ;
                            ROM0_b9     <=  ROM0_arr[12][9]  ;
                            ROM0_b10    <=  ROM0_arr[12][10] ;
                            ROM0_b11    <=  ROM0_arr[12][11] ;
                            ROM0_b12    <=  ROM0_arr[12][12] ;
                            ROM0_b13    <=  ROM0_arr[12][13] ;
                            ROM0_b14    <=  ROM0_arr[12][14] ;
                            ROM0_b15    <=  ROM0_arr[12][15] ;
                        end
                    4'd13:
                        begin
                            ROM0_b0     <=  ROM0_arr[13][0]  ;
                            ROM0_b1     <=  ROM0_arr[13][1]  ;
                            ROM0_b2     <=  ROM0_arr[13][2]  ;
                            ROM0_b3     <=  ROM0_arr[13][3]  ;
                            ROM0_b4     <=  ROM0_arr[13][4]  ;
                            ROM0_b5     <=  ROM0_arr[13][5]  ;
                            ROM0_b6     <=  ROM0_arr[13][6]  ;
                            ROM0_b7     <=  ROM0_arr[13][7]  ;
                            ROM0_b8     <=  ROM0_arr[13][8]  ;
                            ROM0_b9     <=  ROM0_arr[13][9]  ;
                            ROM0_b10    <=  ROM0_arr[13][10] ;
                            ROM0_b11    <=  ROM0_arr[13][11] ;
                            ROM0_b12    <=  ROM0_arr[13][12] ;
                            ROM0_b13    <=  ROM0_arr[13][13] ;
                            ROM0_b14    <=  ROM0_arr[13][14] ;
                            ROM0_b15    <=  ROM0_arr[13][15] ;
                        end
                    4'd14:
                        begin
                            ROM0_b0     <=  ROM0_arr[14][0]  ;
                            ROM0_b1     <=  ROM0_arr[14][1]  ;
                            ROM0_b2     <=  ROM0_arr[14][2]  ;
                            ROM0_b3     <=  ROM0_arr[14][3]  ;
                            ROM0_b4     <=  ROM0_arr[14][4]  ;
                            ROM0_b5     <=  ROM0_arr[14][5]  ;
                            ROM0_b6     <=  ROM0_arr[14][6]  ;
                            ROM0_b7     <=  ROM0_arr[14][7]  ;
                            ROM0_b8     <=  ROM0_arr[14][8]  ;
                            ROM0_b9     <=  ROM0_arr[14][9]  ;
                            ROM0_b10    <=  ROM0_arr[14][10] ;
                            ROM0_b11    <=  ROM0_arr[14][11] ;
                            ROM0_b12    <=  ROM0_arr[14][12] ;
                            ROM0_b13    <=  ROM0_arr[14][13] ;
                            ROM0_b14    <=  ROM0_arr[14][14] ;
                            ROM0_b15    <=  ROM0_arr[14][15] ;
                        end
                    4'd15:
                        begin
                            ROM0_b0     <=  ROM0_arr[15][0]  ;
                            ROM0_b1     <=  ROM0_arr[15][1]  ;
                            ROM0_b2     <=  ROM0_arr[15][2]  ;
                            ROM0_b3     <=  ROM0_arr[15][3]  ;
                            ROM0_b4     <=  ROM0_arr[15][4]  ;
                            ROM0_b5     <=  ROM0_arr[15][5]  ;
                            ROM0_b6     <=  ROM0_arr[15][6]  ;
                            ROM0_b7     <=  ROM0_arr[15][7]  ;
                            ROM0_b8     <=  ROM0_arr[15][8]  ;
                            ROM0_b9     <=  ROM0_arr[15][9]  ;
                            ROM0_b10    <=  ROM0_arr[15][10] ;
                            ROM0_b11    <=  ROM0_arr[15][11] ;
                            ROM0_b12    <=  ROM0_arr[15][12] ;
                            ROM0_b13    <=  ROM0_arr[15][13] ;
                            ROM0_b14    <=  ROM0_arr[15][14] ;
                            ROM0_b15    <=  ROM0_arr[15][15] ;
                        end
                endcase
            end
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM1_b0     <= 64'd0    ;
            ROM1_b1     <= 64'd0    ;
            ROM1_b2     <= 64'd0    ;
            ROM1_b3     <= 64'd0    ;
            ROM1_b4     <= 64'd0    ;
            ROM1_b5     <= 64'd0    ;
            ROM1_b6     <= 64'd0    ;
            ROM1_b7     <= 64'd0    ;
            ROM1_b8     <= 64'd0    ;
            ROM1_b9     <= 64'd0    ;
            ROM1_b10    <= 64'd0    ;
            ROM1_b11    <= 64'd0    ;
            ROM1_b12    <= 64'd0    ; 
            ROM1_b13    <= 64'd0    ;
            ROM1_b14    <= 64'd0    ; 
            ROM1_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (MA1)
                    4'd0:
                        begin
                            ROM1_b0     <=  ROM1_arr[0][0]  ;
                            ROM1_b1     <=  ROM1_arr[0][1]  ;
                            ROM1_b2     <=  ROM1_arr[0][2]  ;
                            ROM1_b3     <=  ROM1_arr[0][3]  ;
                            ROM1_b4     <=  ROM1_arr[0][4]  ;
                            ROM1_b5     <=  ROM1_arr[0][5]  ;
                            ROM1_b6     <=  ROM1_arr[0][6]  ;
                            ROM1_b7     <=  ROM1_arr[0][7]  ;
                            ROM1_b8     <=  ROM1_arr[0][8]  ;
                            ROM1_b9     <=  ROM1_arr[0][9]  ;
                            ROM1_b10    <=  ROM1_arr[0][10] ;
                            ROM1_b11    <=  ROM1_arr[0][11] ;
                            ROM1_b12    <=  ROM1_arr[0][12] ;
                            ROM1_b13    <=  ROM1_arr[0][13] ;
                            ROM1_b14    <=  ROM1_arr[0][14] ;
                            ROM1_b15    <=  ROM1_arr[0][15] ;
                        end
                    4'd1:
                        begin
                            ROM1_b0     <=  ROM1_arr[1][0]  ;
                            ROM1_b1     <=  ROM1_arr[1][1]  ;
                            ROM1_b2     <=  ROM1_arr[1][2]  ;
                            ROM1_b3     <=  ROM1_arr[1][3]  ;
                            ROM1_b4     <=  ROM1_arr[1][4]  ;
                            ROM1_b5     <=  ROM1_arr[1][5]  ;
                            ROM1_b6     <=  ROM1_arr[1][6]  ;
                            ROM1_b7     <=  ROM1_arr[1][7]  ;
                            ROM1_b8     <=  ROM1_arr[1][8]  ;
                            ROM1_b9     <=  ROM1_arr[1][9]  ;
                            ROM1_b10    <=  ROM1_arr[1][10] ;
                            ROM1_b11    <=  ROM1_arr[1][11] ;
                            ROM1_b12    <=  ROM1_arr[1][12] ;
                            ROM1_b13    <=  ROM1_arr[1][13] ;
                            ROM1_b14    <=  ROM1_arr[1][14] ;
                            ROM1_b15    <=  ROM1_arr[1][15] ;
                        end
                    4'd2:
                        begin
                            ROM1_b0     <=  ROM1_arr[2][0]  ;
                            ROM1_b1     <=  ROM1_arr[2][1]  ;
                            ROM1_b2     <=  ROM1_arr[2][2]  ;
                            ROM1_b3     <=  ROM1_arr[2][3]  ;
                            ROM1_b4     <=  ROM1_arr[2][4]  ;
                            ROM1_b5     <=  ROM1_arr[2][5]  ;
                            ROM1_b6     <=  ROM1_arr[2][6]  ;
                            ROM1_b7     <=  ROM1_arr[2][7]  ;
                            ROM1_b8     <=  ROM1_arr[2][8]  ;
                            ROM1_b9     <=  ROM1_arr[2][9]  ;
                            ROM1_b10    <=  ROM1_arr[2][10] ;
                            ROM1_b11    <=  ROM1_arr[2][11] ;
                            ROM1_b12    <=  ROM1_arr[2][12] ;
                            ROM1_b13    <=  ROM1_arr[2][13] ;
                            ROM1_b14    <=  ROM1_arr[2][14] ;
                            ROM1_b15    <=  ROM1_arr[2][15] ;
                        end
                    4'd3:
                        begin
                            ROM1_b0     <=  ROM1_arr[3][0]  ;
                            ROM1_b1     <=  ROM1_arr[3][1]  ;
                            ROM1_b2     <=  ROM1_arr[3][2]  ;
                            ROM1_b3     <=  ROM1_arr[3][3]  ;
                            ROM1_b4     <=  ROM1_arr[3][4]  ;
                            ROM1_b5     <=  ROM1_arr[3][5]  ;
                            ROM1_b6     <=  ROM1_arr[3][6]  ;
                            ROM1_b7     <=  ROM1_arr[3][7]  ;
                            ROM1_b8     <=  ROM1_arr[3][8]  ;
                            ROM1_b9     <=  ROM1_arr[3][9]  ;
                            ROM1_b10    <=  ROM1_arr[3][10] ;
                            ROM1_b11    <=  ROM1_arr[3][11] ;
                            ROM1_b12    <=  ROM1_arr[3][12] ;
                            ROM1_b13    <=  ROM1_arr[3][13] ;
                            ROM1_b14    <=  ROM1_arr[3][14] ;
                            ROM1_b15    <=  ROM1_arr[3][15] ;
                        end
                    4'd4:
                        begin
                            ROM1_b0     <=  ROM1_arr[4][0]  ;
                            ROM1_b1     <=  ROM1_arr[4][1]  ;
                            ROM1_b2     <=  ROM1_arr[4][2]  ;
                            ROM1_b3     <=  ROM1_arr[4][3]  ;
                            ROM1_b4     <=  ROM1_arr[4][4]  ;
                            ROM1_b5     <=  ROM1_arr[4][5]  ;
                            ROM1_b6     <=  ROM1_arr[4][6]  ;
                            ROM1_b7     <=  ROM1_arr[4][7]  ;
                            ROM1_b8     <=  ROM1_arr[4][8]  ;
                            ROM1_b9     <=  ROM1_arr[4][9]  ;
                            ROM1_b10    <=  ROM1_arr[4][10] ;
                            ROM1_b11    <=  ROM1_arr[4][11] ;
                            ROM1_b12    <=  ROM1_arr[4][12] ;
                            ROM1_b13    <=  ROM1_arr[4][13] ;
                            ROM1_b14    <=  ROM1_arr[4][14] ;
                            ROM1_b15    <=  ROM1_arr[4][15] ;
                        end
                    4'd5:
                        begin
                            ROM1_b0     <=  ROM1_arr[5][0]  ;
                            ROM1_b1     <=  ROM1_arr[5][1]  ;
                            ROM1_b2     <=  ROM1_arr[5][2]  ;
                            ROM1_b3     <=  ROM1_arr[5][3]  ;
                            ROM1_b4     <=  ROM1_arr[5][4]  ;
                            ROM1_b5     <=  ROM1_arr[5][5]  ;
                            ROM1_b6     <=  ROM1_arr[5][6]  ;
                            ROM1_b7     <=  ROM1_arr[5][7]  ;
                            ROM1_b8     <=  ROM1_arr[5][8]  ;
                            ROM1_b9     <=  ROM1_arr[5][9]  ;
                            ROM1_b10    <=  ROM1_arr[5][10] ;
                            ROM1_b11    <=  ROM1_arr[5][11] ;
                            ROM1_b12    <=  ROM1_arr[5][12] ;
                            ROM1_b13    <=  ROM1_arr[5][13] ;
                            ROM1_b14    <=  ROM1_arr[5][14] ;
                            ROM1_b15    <=  ROM1_arr[5][15] ;
                        end
                    4'd6:
                        begin
                            ROM1_b0     <=  ROM1_arr[6][0]  ;
                            ROM1_b1     <=  ROM1_arr[6][1]  ;
                            ROM1_b2     <=  ROM1_arr[6][2]  ;
                            ROM1_b3     <=  ROM1_arr[6][3]  ;
                            ROM1_b4     <=  ROM1_arr[6][4]  ;
                            ROM1_b5     <=  ROM1_arr[6][5]  ;
                            ROM1_b6     <=  ROM1_arr[6][6]  ;
                            ROM1_b7     <=  ROM1_arr[6][7]  ;
                            ROM1_b8     <=  ROM1_arr[6][8]  ;
                            ROM1_b9     <=  ROM1_arr[6][9]  ;
                            ROM1_b10    <=  ROM1_arr[6][10] ;
                            ROM1_b11    <=  ROM1_arr[6][11] ;
                            ROM1_b12    <=  ROM1_arr[6][12] ;
                            ROM1_b13    <=  ROM1_arr[6][13] ;
                            ROM1_b14    <=  ROM1_arr[6][14] ;
                            ROM1_b15    <=  ROM1_arr[6][15] ;
                        end
                    4'd7:
                        begin
                            ROM1_b0     <=  ROM1_arr[7][0]  ;
                            ROM1_b1     <=  ROM1_arr[7][1]  ;
                            ROM1_b2     <=  ROM1_arr[7][2]  ;
                            ROM1_b3     <=  ROM1_arr[7][3]  ;
                            ROM1_b4     <=  ROM1_arr[7][4]  ;
                            ROM1_b5     <=  ROM1_arr[7][5]  ;
                            ROM1_b6     <=  ROM1_arr[7][6]  ;
                            ROM1_b7     <=  ROM1_arr[7][7]  ;
                            ROM1_b8     <=  ROM1_arr[7][8]  ;
                            ROM1_b9     <=  ROM1_arr[7][9]  ;
                            ROM1_b10    <=  ROM1_arr[7][10] ;
                            ROM1_b11    <=  ROM1_arr[7][11] ;
                            ROM1_b12    <=  ROM1_arr[7][12] ;
                            ROM1_b13    <=  ROM1_arr[7][13] ;
                            ROM1_b14    <=  ROM1_arr[7][14] ;
                            ROM1_b15    <=  ROM1_arr[7][15] ;
                        end
                    4'd8:
                        begin
                            ROM1_b0     <=  ROM1_arr[8][0]  ;
                            ROM1_b1     <=  ROM1_arr[8][1]  ;
                            ROM1_b2     <=  ROM1_arr[8][2]  ;
                            ROM1_b3     <=  ROM1_arr[8][3]  ;
                            ROM1_b4     <=  ROM1_arr[8][4]  ;
                            ROM1_b5     <=  ROM1_arr[8][5]  ;
                            ROM1_b6     <=  ROM1_arr[8][6]  ;
                            ROM1_b7     <=  ROM1_arr[8][7]  ;
                            ROM1_b8     <=  ROM1_arr[8][8]  ;
                            ROM1_b9     <=  ROM1_arr[8][9]  ;
                            ROM1_b10    <=  ROM1_arr[8][10] ;
                            ROM1_b11    <=  ROM1_arr[8][11] ;
                            ROM1_b12    <=  ROM1_arr[8][12] ;
                            ROM1_b13    <=  ROM1_arr[8][13] ;
                            ROM1_b14    <=  ROM1_arr[8][14] ;
                            ROM1_b15    <=  ROM1_arr[8][15] ;
                        end
                    4'd9:
                        begin
                            ROM1_b0     <=  ROM1_arr[9][0]  ;
                            ROM1_b1     <=  ROM1_arr[9][1]  ;
                            ROM1_b2     <=  ROM1_arr[9][2]  ;
                            ROM1_b3     <=  ROM1_arr[9][3]  ;
                            ROM1_b4     <=  ROM1_arr[9][4]  ;
                            ROM1_b5     <=  ROM1_arr[9][5]  ;
                            ROM1_b6     <=  ROM1_arr[9][6]  ;
                            ROM1_b7     <=  ROM1_arr[9][7]  ;
                            ROM1_b8     <=  ROM1_arr[9][8]  ;
                            ROM1_b9     <=  ROM1_arr[9][9]  ;
                            ROM1_b10    <=  ROM1_arr[9][10] ;
                            ROM1_b11    <=  ROM1_arr[9][11] ;
                            ROM1_b12    <=  ROM1_arr[9][12] ;
                            ROM1_b13    <=  ROM1_arr[9][13] ;
                            ROM1_b14    <=  ROM1_arr[9][14] ;
                            ROM1_b15    <=  ROM1_arr[9][15] ;
                        end
                    4'd10:
                        begin
                            ROM1_b0     <=  ROM1_arr[10][0]  ;
                            ROM1_b1     <=  ROM1_arr[10][1]  ;
                            ROM1_b2     <=  ROM1_arr[10][2]  ;
                            ROM1_b3     <=  ROM1_arr[10][3]  ;
                            ROM1_b4     <=  ROM1_arr[10][4]  ;
                            ROM1_b5     <=  ROM1_arr[10][5]  ;
                            ROM1_b6     <=  ROM1_arr[10][6]  ;
                            ROM1_b7     <=  ROM1_arr[10][7]  ;
                            ROM1_b8     <=  ROM1_arr[10][8]  ;
                            ROM1_b9     <=  ROM1_arr[10][9]  ;
                            ROM1_b10    <=  ROM1_arr[10][10] ;
                            ROM1_b11    <=  ROM1_arr[10][11] ;
                            ROM1_b12    <=  ROM1_arr[10][12] ;
                            ROM1_b13    <=  ROM1_arr[10][13] ;
                            ROM1_b14    <=  ROM1_arr[10][14] ;
                            ROM1_b15    <=  ROM1_arr[10][15] ;
                        end
                    4'd11:
                        begin
                            ROM1_b0     <=  ROM1_arr[11][0]  ;
                            ROM1_b1     <=  ROM1_arr[11][1]  ;
                            ROM1_b2     <=  ROM1_arr[11][2]  ;
                            ROM1_b3     <=  ROM1_arr[11][3]  ;
                            ROM1_b4     <=  ROM1_arr[11][4]  ;
                            ROM1_b5     <=  ROM1_arr[11][5]  ;
                            ROM1_b6     <=  ROM1_arr[11][6]  ;
                            ROM1_b7     <=  ROM1_arr[11][7]  ;
                            ROM1_b8     <=  ROM1_arr[11][8]  ;
                            ROM1_b9     <=  ROM1_arr[11][9]  ;
                            ROM1_b10    <=  ROM1_arr[11][10] ;
                            ROM1_b11    <=  ROM1_arr[11][11] ;
                            ROM1_b12    <=  ROM1_arr[11][12] ;
                            ROM1_b13    <=  ROM1_arr[11][13] ;
                            ROM1_b14    <=  ROM1_arr[11][14] ;
                            ROM1_b15    <=  ROM1_arr[11][15] ;
                        end
                    4'd12:
                        begin
                            ROM1_b0     <=  ROM1_arr[12][0]  ;
                            ROM1_b1     <=  ROM1_arr[12][1]  ;
                            ROM1_b2     <=  ROM1_arr[12][2]  ;
                            ROM1_b3     <=  ROM1_arr[12][3]  ;
                            ROM1_b4     <=  ROM1_arr[12][4]  ;
                            ROM1_b5     <=  ROM1_arr[12][5]  ;
                            ROM1_b6     <=  ROM1_arr[12][6]  ;
                            ROM1_b7     <=  ROM1_arr[12][7]  ;
                            ROM1_b8     <=  ROM1_arr[12][8]  ;
                            ROM1_b9     <=  ROM1_arr[12][9]  ;
                            ROM1_b10    <=  ROM1_arr[12][10] ;
                            ROM1_b11    <=  ROM1_arr[12][11] ;
                            ROM1_b12    <=  ROM1_arr[12][12] ;
                            ROM1_b13    <=  ROM1_arr[12][13] ;
                            ROM1_b14    <=  ROM1_arr[12][14] ;
                            ROM1_b15    <=  ROM1_arr[12][15] ;
                        end
                    4'd13:
                        begin
                            ROM1_b0     <=  ROM1_arr[13][0]  ;
                            ROM1_b1     <=  ROM1_arr[13][1]  ;
                            ROM1_b2     <=  ROM1_arr[13][2]  ;
                            ROM1_b3     <=  ROM1_arr[13][3]  ;
                            ROM1_b4     <=  ROM1_arr[13][4]  ;
                            ROM1_b5     <=  ROM1_arr[13][5]  ;
                            ROM1_b6     <=  ROM1_arr[13][6]  ;
                            ROM1_b7     <=  ROM1_arr[13][7]  ;
                            ROM1_b8     <=  ROM1_arr[13][8]  ;
                            ROM1_b9     <=  ROM1_arr[13][9]  ;
                            ROM1_b10    <=  ROM1_arr[13][10] ;
                            ROM1_b11    <=  ROM1_arr[13][11] ;
                            ROM1_b12    <=  ROM1_arr[13][12] ;
                            ROM1_b13    <=  ROM1_arr[13][13] ;
                            ROM1_b14    <=  ROM1_arr[13][14] ;
                            ROM1_b15    <=  ROM1_arr[13][15] ;
                        end
                    4'd14:
                        begin
                            ROM1_b0     <=  ROM1_arr[14][0]  ;
                            ROM1_b1     <=  ROM1_arr[14][1]  ;
                            ROM1_b2     <=  ROM1_arr[14][2]  ;
                            ROM1_b3     <=  ROM1_arr[14][3]  ;
                            ROM1_b4     <=  ROM1_arr[14][4]  ;
                            ROM1_b5     <=  ROM1_arr[14][5]  ;
                            ROM1_b6     <=  ROM1_arr[14][6]  ;
                            ROM1_b7     <=  ROM1_arr[14][7]  ;
                            ROM1_b8     <=  ROM1_arr[14][8]  ;
                            ROM1_b9     <=  ROM1_arr[14][9]  ;
                            ROM1_b10    <=  ROM1_arr[14][10] ;
                            ROM1_b11    <=  ROM1_arr[14][11] ;
                            ROM1_b12    <=  ROM1_arr[14][12] ;
                            ROM1_b13    <=  ROM1_arr[14][13] ;
                            ROM1_b14    <=  ROM1_arr[14][14] ;
                            ROM1_b15    <=  ROM1_arr[14][15] ;
                        end
                    4'd15:
                        begin
                            ROM1_b0     <=  ROM1_arr[15][0]  ;
                            ROM1_b1     <=  ROM1_arr[15][1]  ;
                            ROM1_b2     <=  ROM1_arr[15][2]  ;
                            ROM1_b3     <=  ROM1_arr[15][3]  ;
                            ROM1_b4     <=  ROM1_arr[15][4]  ;
                            ROM1_b5     <=  ROM1_arr[15][5]  ;
                            ROM1_b6     <=  ROM1_arr[15][6]  ;
                            ROM1_b7     <=  ROM1_arr[15][7]  ;
                            ROM1_b8     <=  ROM1_arr[15][8]  ;
                            ROM1_b9     <=  ROM1_arr[15][9]  ;
                            ROM1_b10    <=  ROM1_arr[15][10] ;
                            ROM1_b11    <=  ROM1_arr[15][11] ;
                            ROM1_b12    <=  ROM1_arr[15][12] ;
                            ROM1_b13    <=  ROM1_arr[15][13] ;
                            ROM1_b14    <=  ROM1_arr[15][14] ;
                            ROM1_b15    <=  ROM1_arr[15][15] ;
                        end
                endcase
            end
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM2_b0     <= 64'd0    ;
            ROM2_b1     <= 64'd0    ;
            ROM2_b2     <= 64'd0    ;
            ROM2_b3     <= 64'd0    ;
            ROM2_b4     <= 64'd0    ;
            ROM2_b5     <= 64'd0    ;
            ROM2_b6     <= 64'd0    ;
            ROM2_b7     <= 64'd0    ;
            ROM2_b8     <= 64'd0    ;
            ROM2_b9     <= 64'd0    ;
            ROM2_b10    <= 64'd0    ;
            ROM2_b11    <= 64'd0    ;
            ROM2_b12    <= 64'd0    ; 
            ROM2_b13    <= 64'd0    ;
            ROM2_b14    <= 64'd0    ; 
            ROM2_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (MA2)
                    4'd0:
                        begin
                            ROM2_b0     <=  ROM2_arr[0][0]  ;
                            ROM2_b1     <=  ROM2_arr[0][1]  ;
                            ROM2_b2     <=  ROM2_arr[0][2]  ;
                            ROM2_b3     <=  ROM2_arr[0][3]  ;
                            ROM2_b4     <=  ROM2_arr[0][4]  ;
                            ROM2_b5     <=  ROM2_arr[0][5]  ;
                            ROM2_b6     <=  ROM2_arr[0][6]  ;
                            ROM2_b7     <=  ROM2_arr[0][7]  ;
                            ROM2_b8     <=  ROM2_arr[0][8]  ;
                            ROM2_b9     <=  ROM2_arr[0][9]  ;
                            ROM2_b10    <=  ROM2_arr[0][10] ;
                            ROM2_b11    <=  ROM2_arr[0][11] ;
                            ROM2_b12    <=  ROM2_arr[0][12] ;
                            ROM2_b13    <=  ROM2_arr[0][13] ;
                            ROM2_b14    <=  ROM2_arr[0][14] ;
                            ROM2_b15    <=  ROM2_arr[0][15] ;
                        end
                    4'd1:
                        begin
                            ROM2_b0     <=  ROM2_arr[1][0]  ;
                            ROM2_b1     <=  ROM2_arr[1][1]  ;
                            ROM2_b2     <=  ROM2_arr[1][2]  ;
                            ROM2_b3     <=  ROM2_arr[1][3]  ;
                            ROM2_b4     <=  ROM2_arr[1][4]  ;
                            ROM2_b5     <=  ROM2_arr[1][5]  ;
                            ROM2_b6     <=  ROM2_arr[1][6]  ;
                            ROM2_b7     <=  ROM2_arr[1][7]  ;
                            ROM2_b8     <=  ROM2_arr[1][8]  ;
                            ROM2_b9     <=  ROM2_arr[1][9]  ;
                            ROM2_b10    <=  ROM2_arr[1][10] ;
                            ROM2_b11    <=  ROM2_arr[1][11] ;
                            ROM2_b12    <=  ROM2_arr[1][12] ;
                            ROM2_b13    <=  ROM2_arr[1][13] ;
                            ROM2_b14    <=  ROM2_arr[1][14] ;
                            ROM2_b15    <=  ROM2_arr[1][15] ;
                        end
                    4'd2:
                        begin
                            ROM2_b0     <=  ROM2_arr[2][0]  ;
                            ROM2_b1     <=  ROM2_arr[2][1]  ;
                            ROM2_b2     <=  ROM2_arr[2][2]  ;
                            ROM2_b3     <=  ROM2_arr[2][3]  ;
                            ROM2_b4     <=  ROM2_arr[2][4]  ;
                            ROM2_b5     <=  ROM2_arr[2][5]  ;
                            ROM2_b6     <=  ROM2_arr[2][6]  ;
                            ROM2_b7     <=  ROM2_arr[2][7]  ;
                            ROM2_b8     <=  ROM2_arr[2][8]  ;
                            ROM2_b9     <=  ROM2_arr[2][9]  ;
                            ROM2_b10    <=  ROM2_arr[2][10] ;
                            ROM2_b11    <=  ROM2_arr[2][11] ;
                            ROM2_b12    <=  ROM2_arr[2][12] ;
                            ROM2_b13    <=  ROM2_arr[2][13] ;
                            ROM2_b14    <=  ROM2_arr[2][14] ;
                            ROM2_b15    <=  ROM2_arr[2][15] ;
                        end
                    4'd3:
                        begin
                            ROM2_b0     <=  ROM2_arr[3][0]  ;
                            ROM2_b1     <=  ROM2_arr[3][1]  ;
                            ROM2_b2     <=  ROM2_arr[3][2]  ;
                            ROM2_b3     <=  ROM2_arr[3][3]  ;
                            ROM2_b4     <=  ROM2_arr[3][4]  ;
                            ROM2_b5     <=  ROM2_arr[3][5]  ;
                            ROM2_b6     <=  ROM2_arr[3][6]  ;
                            ROM2_b7     <=  ROM2_arr[3][7]  ;
                            ROM2_b8     <=  ROM2_arr[3][8]  ;
                            ROM2_b9     <=  ROM2_arr[3][9]  ;
                            ROM2_b10    <=  ROM2_arr[3][10] ;
                            ROM2_b11    <=  ROM2_arr[3][11] ;
                            ROM2_b12    <=  ROM2_arr[3][12] ;
                            ROM2_b13    <=  ROM2_arr[3][13] ;
                            ROM2_b14    <=  ROM2_arr[3][14] ;
                            ROM2_b15    <=  ROM2_arr[3][15] ;
                        end
                    4'd4:
                        begin
                            ROM2_b0     <=  ROM2_arr[4][0]  ;
                            ROM2_b1     <=  ROM2_arr[4][1]  ;
                            ROM2_b2     <=  ROM2_arr[4][2]  ;
                            ROM2_b3     <=  ROM2_arr[4][3]  ;
                            ROM2_b4     <=  ROM2_arr[4][4]  ;
                            ROM2_b5     <=  ROM2_arr[4][5]  ;
                            ROM2_b6     <=  ROM2_arr[4][6]  ;
                            ROM2_b7     <=  ROM2_arr[4][7]  ;
                            ROM2_b8     <=  ROM2_arr[4][8]  ;
                            ROM2_b9     <=  ROM2_arr[4][9]  ;
                            ROM2_b10    <=  ROM2_arr[4][10] ;
                            ROM2_b11    <=  ROM2_arr[4][11] ;
                            ROM2_b12    <=  ROM2_arr[4][12] ;
                            ROM2_b13    <=  ROM2_arr[4][13] ;
                            ROM2_b14    <=  ROM2_arr[4][14] ;
                            ROM2_b15    <=  ROM2_arr[4][15] ;
                        end
                    4'd5:
                        begin
                            ROM2_b0     <=  ROM2_arr[5][0]  ;
                            ROM2_b1     <=  ROM2_arr[5][1]  ;
                            ROM2_b2     <=  ROM2_arr[5][2]  ;
                            ROM2_b3     <=  ROM2_arr[5][3]  ;
                            ROM2_b4     <=  ROM2_arr[5][4]  ;
                            ROM2_b5     <=  ROM2_arr[5][5]  ;
                            ROM2_b6     <=  ROM2_arr[5][6]  ;
                            ROM2_b7     <=  ROM2_arr[5][7]  ;
                            ROM2_b8     <=  ROM2_arr[5][8]  ;
                            ROM2_b9     <=  ROM2_arr[5][9]  ;
                            ROM2_b10    <=  ROM2_arr[5][10] ;
                            ROM2_b11    <=  ROM2_arr[5][11] ;
                            ROM2_b12    <=  ROM2_arr[5][12] ;
                            ROM2_b13    <=  ROM2_arr[5][13] ;
                            ROM2_b14    <=  ROM2_arr[5][14] ;
                            ROM2_b15    <=  ROM2_arr[5][15] ;
                        end
                    4'd6:
                        begin
                            ROM2_b0     <=  ROM2_arr[6][0]  ;
                            ROM2_b1     <=  ROM2_arr[6][1]  ;
                            ROM2_b2     <=  ROM2_arr[6][2]  ;
                            ROM2_b3     <=  ROM2_arr[6][3]  ;
                            ROM2_b4     <=  ROM2_arr[6][4]  ;
                            ROM2_b5     <=  ROM2_arr[6][5]  ;
                            ROM2_b6     <=  ROM2_arr[6][6]  ;
                            ROM2_b7     <=  ROM2_arr[6][7]  ;
                            ROM2_b8     <=  ROM2_arr[6][8]  ;
                            ROM2_b9     <=  ROM2_arr[6][9]  ;
                            ROM2_b10    <=  ROM2_arr[6][10] ;
                            ROM2_b11    <=  ROM2_arr[6][11] ;
                            ROM2_b12    <=  ROM2_arr[6][12] ;
                            ROM2_b13    <=  ROM2_arr[6][13] ;
                            ROM2_b14    <=  ROM2_arr[6][14] ;
                            ROM2_b15    <=  ROM2_arr[6][15] ;
                        end
                    4'd7:
                        begin
                            ROM2_b0     <=  ROM2_arr[7][0]  ;
                            ROM2_b1     <=  ROM2_arr[7][1]  ;
                            ROM2_b2     <=  ROM2_arr[7][2]  ;
                            ROM2_b3     <=  ROM2_arr[7][3]  ;
                            ROM2_b4     <=  ROM2_arr[7][4]  ;
                            ROM2_b5     <=  ROM2_arr[7][5]  ;
                            ROM2_b6     <=  ROM2_arr[7][6]  ;
                            ROM2_b7     <=  ROM2_arr[7][7]  ;
                            ROM2_b8     <=  ROM2_arr[7][8]  ;
                            ROM2_b9     <=  ROM2_arr[7][9]  ;
                            ROM2_b10    <=  ROM2_arr[7][10] ;
                            ROM2_b11    <=  ROM2_arr[7][11] ;
                            ROM2_b12    <=  ROM2_arr[7][12] ;
                            ROM2_b13    <=  ROM2_arr[7][13] ;
                            ROM2_b14    <=  ROM2_arr[7][14] ;
                            ROM2_b15    <=  ROM2_arr[7][15] ;
                        end
                    4'd8:
                        begin
                            ROM2_b0     <=  ROM2_arr[8][0]  ;
                            ROM2_b1     <=  ROM2_arr[8][1]  ;
                            ROM2_b2     <=  ROM2_arr[8][2]  ;
                            ROM2_b3     <=  ROM2_arr[8][3]  ;
                            ROM2_b4     <=  ROM2_arr[8][4]  ;
                            ROM2_b5     <=  ROM2_arr[8][5]  ;
                            ROM2_b6     <=  ROM2_arr[8][6]  ;
                            ROM2_b7     <=  ROM2_arr[8][7]  ;
                            ROM2_b8     <=  ROM2_arr[8][8]  ;
                            ROM2_b9     <=  ROM2_arr[8][9]  ;
                            ROM2_b10    <=  ROM2_arr[8][10] ;
                            ROM2_b11    <=  ROM2_arr[8][11] ;
                            ROM2_b12    <=  ROM2_arr[8][12] ;
                            ROM2_b13    <=  ROM2_arr[8][13] ;
                            ROM2_b14    <=  ROM2_arr[8][14] ;
                            ROM2_b15    <=  ROM2_arr[8][15] ;
                        end
                    4'd9:
                        begin
                            ROM2_b0     <=  ROM2_arr[9][0]  ;
                            ROM2_b1     <=  ROM2_arr[9][1]  ;
                            ROM2_b2     <=  ROM2_arr[9][2]  ;
                            ROM2_b3     <=  ROM2_arr[9][3]  ;
                            ROM2_b4     <=  ROM2_arr[9][4]  ;
                            ROM2_b5     <=  ROM2_arr[9][5]  ;
                            ROM2_b6     <=  ROM2_arr[9][6]  ;
                            ROM2_b7     <=  ROM2_arr[9][7]  ;
                            ROM2_b8     <=  ROM2_arr[9][8]  ;
                            ROM2_b9     <=  ROM2_arr[9][9]  ;
                            ROM2_b10    <=  ROM2_arr[9][10] ;
                            ROM2_b11    <=  ROM2_arr[9][11] ;
                            ROM2_b12    <=  ROM2_arr[9][12] ;
                            ROM2_b13    <=  ROM2_arr[9][13] ;
                            ROM2_b14    <=  ROM2_arr[9][14] ;
                            ROM2_b15    <=  ROM2_arr[9][15] ;
                        end
                    4'd10:
                        begin
                            ROM2_b0     <=  ROM2_arr[10][0]  ;
                            ROM2_b1     <=  ROM2_arr[10][1]  ;
                            ROM2_b2     <=  ROM2_arr[10][2]  ;
                            ROM2_b3     <=  ROM2_arr[10][3]  ;
                            ROM2_b4     <=  ROM2_arr[10][4]  ;
                            ROM2_b5     <=  ROM2_arr[10][5]  ;
                            ROM2_b6     <=  ROM2_arr[10][6]  ;
                            ROM2_b7     <=  ROM2_arr[10][7]  ;
                            ROM2_b8     <=  ROM2_arr[10][8]  ;
                            ROM2_b9     <=  ROM2_arr[10][9]  ;
                            ROM2_b10    <=  ROM2_arr[10][10] ;
                            ROM2_b11    <=  ROM2_arr[10][11] ;
                            ROM2_b12    <=  ROM2_arr[10][12] ;
                            ROM2_b13    <=  ROM2_arr[10][13] ;
                            ROM2_b14    <=  ROM2_arr[10][14] ;
                            ROM2_b15    <=  ROM2_arr[10][15] ;
                        end
                    4'd11:
                        begin
                            ROM2_b0     <=  ROM2_arr[11][0]  ;
                            ROM2_b1     <=  ROM2_arr[11][1]  ;
                            ROM2_b2     <=  ROM2_arr[11][2]  ;
                            ROM2_b3     <=  ROM2_arr[11][3]  ;
                            ROM2_b4     <=  ROM2_arr[11][4]  ;
                            ROM2_b5     <=  ROM2_arr[11][5]  ;
                            ROM2_b6     <=  ROM2_arr[11][6]  ;
                            ROM2_b7     <=  ROM2_arr[11][7]  ;
                            ROM2_b8     <=  ROM2_arr[11][8]  ;
                            ROM2_b9     <=  ROM2_arr[11][9]  ;
                            ROM2_b10    <=  ROM2_arr[11][10] ;
                            ROM2_b11    <=  ROM2_arr[11][11] ;
                            ROM2_b12    <=  ROM2_arr[11][12] ;
                            ROM2_b13    <=  ROM2_arr[11][13] ;
                            ROM2_b14    <=  ROM2_arr[11][14] ;
                            ROM2_b15    <=  ROM2_arr[11][15] ;
                        end
                    4'd12:
                        begin
                            ROM2_b0     <=  ROM2_arr[12][0]  ;
                            ROM2_b1     <=  ROM2_arr[12][1]  ;
                            ROM2_b2     <=  ROM2_arr[12][2]  ;
                            ROM2_b3     <=  ROM2_arr[12][3]  ;
                            ROM2_b4     <=  ROM2_arr[12][4]  ;
                            ROM2_b5     <=  ROM2_arr[12][5]  ;
                            ROM2_b6     <=  ROM2_arr[12][6]  ;
                            ROM2_b7     <=  ROM2_arr[12][7]  ;
                            ROM2_b8     <=  ROM2_arr[12][8]  ;
                            ROM2_b9     <=  ROM2_arr[12][9]  ;
                            ROM2_b10    <=  ROM2_arr[12][10] ;
                            ROM2_b11    <=  ROM2_arr[12][11] ;
                            ROM2_b12    <=  ROM2_arr[12][12] ;
                            ROM2_b13    <=  ROM2_arr[12][13] ;
                            ROM2_b14    <=  ROM2_arr[12][14] ;
                            ROM2_b15    <=  ROM2_arr[12][15] ;
                        end
                    4'd13:
                        begin
                            ROM2_b0     <=  ROM2_arr[13][0]  ;
                            ROM2_b1     <=  ROM2_arr[13][1]  ;
                            ROM2_b2     <=  ROM2_arr[13][2]  ;
                            ROM2_b3     <=  ROM2_arr[13][3]  ;
                            ROM2_b4     <=  ROM2_arr[13][4]  ;
                            ROM2_b5     <=  ROM2_arr[13][5]  ;
                            ROM2_b6     <=  ROM2_arr[13][6]  ;
                            ROM2_b7     <=  ROM2_arr[13][7]  ;
                            ROM2_b8     <=  ROM2_arr[13][8]  ;
                            ROM2_b9     <=  ROM2_arr[13][9]  ;
                            ROM2_b10    <=  ROM2_arr[13][10] ;
                            ROM2_b11    <=  ROM2_arr[13][11] ;
                            ROM2_b12    <=  ROM2_arr[13][12] ;
                            ROM2_b13    <=  ROM2_arr[13][13] ;
                            ROM2_b14    <=  ROM2_arr[13][14] ;
                            ROM2_b15    <=  ROM2_arr[13][15] ;
                        end
                    4'd14:
                        begin
                            ROM2_b0     <=  ROM2_arr[14][0]  ;
                            ROM2_b1     <=  ROM2_arr[14][1]  ;
                            ROM2_b2     <=  ROM2_arr[14][2]  ;
                            ROM2_b3     <=  ROM2_arr[14][3]  ;
                            ROM2_b4     <=  ROM2_arr[14][4]  ;
                            ROM2_b5     <=  ROM2_arr[14][5]  ;
                            ROM2_b6     <=  ROM2_arr[14][6]  ;
                            ROM2_b7     <=  ROM2_arr[14][7]  ;
                            ROM2_b8     <=  ROM2_arr[14][8]  ;
                            ROM2_b9     <=  ROM2_arr[14][9]  ;
                            ROM2_b10    <=  ROM2_arr[14][10] ;
                            ROM2_b11    <=  ROM2_arr[14][11] ;
                            ROM2_b12    <=  ROM2_arr[14][12] ;
                            ROM2_b13    <=  ROM2_arr[14][13] ;
                            ROM2_b14    <=  ROM2_arr[14][14] ;
                            ROM2_b15    <=  ROM2_arr[14][15] ;
                        end
                    4'd15:
                        begin
                            ROM2_b0     <=  ROM2_arr[15][0]  ;
                            ROM2_b1     <=  ROM2_arr[15][1]  ;
                            ROM2_b2     <=  ROM2_arr[15][2]  ;
                            ROM2_b3     <=  ROM2_arr[15][3]  ;
                            ROM2_b4     <=  ROM2_arr[15][4]  ;
                            ROM2_b5     <=  ROM2_arr[15][5]  ;
                            ROM2_b6     <=  ROM2_arr[15][6]  ;
                            ROM2_b7     <=  ROM2_arr[15][7]  ;
                            ROM2_b8     <=  ROM2_arr[15][8]  ;
                            ROM2_b9     <=  ROM2_arr[15][9]  ;
                            ROM2_b10    <=  ROM2_arr[15][10] ;
                            ROM2_b11    <=  ROM2_arr[15][11] ;
                            ROM2_b12    <=  ROM2_arr[15][12] ;
                            ROM2_b13    <=  ROM2_arr[15][13] ;
                            ROM2_b14    <=  ROM2_arr[15][14] ;
                            ROM2_b15    <=  ROM2_arr[15][15] ;
                        end
                endcase
            end
        end
    end
endmodule