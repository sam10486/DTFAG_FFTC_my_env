`include "define.v"
module Register_file (
    input clk,
    input rst_n,
    input [`ROMA_width-1:0] MA0,
    input [`ROMA_width-1:0] MA1,
    input [`ROMA_width-1:0] MA2,
    input ROM_CEN,
    input [1:0] FFT_stage_in,

    output reg [`D_width-1:0] ROM0_b0   ,
    output reg [`D_width-1:0] ROM0_b1   ,
    output reg [`D_width-1:0] ROM0_b2   ,
    output reg [`D_width-1:0] ROM0_b3   ,
    output reg [`D_width-1:0] ROM0_b4   ,
    output reg [`D_width-1:0] ROM0_b5   ,
    output reg [`D_width-1:0] ROM0_b6   ,
    output reg [`D_width-1:0] ROM0_b7   ,
    output reg [`D_width-1:0] ROM0_b8   ,
    output reg [`D_width-1:0] ROM0_b9   ,
    output reg [`D_width-1:0] ROM0_b10  ,
    output reg [`D_width-1:0] ROM0_b11  ,
    output reg [`D_width-1:0] ROM0_b12  ,
    output reg [`D_width-1:0] ROM0_b13  ,
    output reg [`D_width-1:0] ROM0_b14  ,
    output reg [`D_width-1:0] ROM0_b15  ,
    // ROM1
    output reg [`D_width-1:0] ROM1_b0   ,
    output reg [`D_width-1:0] ROM1_b1   ,
    output reg [`D_width-1:0] ROM1_b2   ,
    output reg [`D_width-1:0] ROM1_b3   ,
    output reg [`D_width-1:0] ROM1_b4   ,
    output reg [`D_width-1:0] ROM1_b5   ,
    output reg [`D_width-1:0] ROM1_b6   ,
    output reg [`D_width-1:0] ROM1_b7   ,
    output reg [`D_width-1:0] ROM1_b8   ,
    output reg [`D_width-1:0] ROM1_b9   ,
    output reg [`D_width-1:0] ROM1_b10  ,
    output reg [`D_width-1:0] ROM1_b11  ,
    output reg [`D_width-1:0] ROM1_b12  ,
    output reg [`D_width-1:0] ROM1_b13  ,
    output reg [`D_width-1:0] ROM1_b14  ,
    output reg [`D_width-1:0] ROM1_b15  ,
    // ROM2
    output reg [`D_width-1:0] ROM2_b0   ,
    output reg [`D_width-1:0] ROM2_b1   ,
    output reg [`D_width-1:0] ROM2_b2   ,
    output reg [`D_width-1:0] ROM2_b3   ,
    output reg [`D_width-1:0] ROM2_b4   ,
    output reg [`D_width-1:0] ROM2_b5   ,
    output reg [`D_width-1:0] ROM2_b6   ,
    output reg [`D_width-1:0] ROM2_b7   ,
    output reg [`D_width-1:0] ROM2_b8   ,
    output reg [`D_width-1:0] ROM2_b9   ,
    output reg [`D_width-1:0] ROM2_b10  ,
    output reg [`D_width-1:0] ROM2_b11  ,
    output reg [`D_width-1:0] ROM2_b12  ,
    output reg [`D_width-1:0] ROM2_b13  ,
    output reg [`D_width-1:0] ROM2_b14  ,
    output reg [`D_width-1:0] ROM2_b15  
);

    reg [`D_width-1:0] ROM0_st0_arr [0:15][0:15];
    reg [`D_width-1:0] ROM0_st1_arr [0:15][0:15];
    reg [`D_width-1:0] ROM0_st2_arr [0:15][0:15];
    reg [`D_width-1:0] ROM0_st3_arr [0:15];
    reg [`D_width-1:0] ROM1_arr [0:15][0:15];
    reg [`D_width-1:0] ROM2_arr [0:15][0:15];
    
    always@( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            // ROM0 init
            ROM0_st0_arr[0][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[0][1] <= 64'd10793526415136183099;
            ROM0_st0_arr[0][2] <= 64'd13209821187581267427;
            ROM0_st0_arr[0][3] <= 64'd264562574883826952;
            ROM0_st0_arr[0][4] <= 64'd16659427319513139460;
            ROM0_st0_arr[0][5] <= 64'd17552852175845899994;
            ROM0_st0_arr[0][6] <= 64'd14396015468671915866;
            ROM0_st0_arr[0][7] <= 64'd5562516121259070392;
            ROM0_st0_arr[0][8] <= 64'd11286921907217085921;
            ROM0_st0_arr[0][9] <= 64'd16754059815999085656;
            ROM0_st0_arr[0][10] <= 64'd15595010439883317588;
            ROM0_st0_arr[0][11] <= 64'd3772231912420796197;
            ROM0_st0_arr[0][12] <= 64'd14367586735222943862;
            ROM0_st0_arr[0][13] <= 64'd14051862940598240066;
            ROM0_st0_arr[0][14] <= 64'd1493072641708298704;
            ROM0_st0_arr[0][15] <= 64'd13344274783299470058;
            ROM0_st0_arr[1][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[1][1] <= 64'd9695816016920606992;
            ROM0_st0_arr[1][2] <= 64'd10296873228810115991;
            ROM0_st0_arr[1][3] <= 64'd50652191562594056;
            ROM0_st0_arr[1][4] <= 64'd16049903969184754810;
            ROM0_st0_arr[1][5] <= 64'd12828076810033474802;
            ROM0_st0_arr[1][6] <= 64'd14977535962704764430;
            ROM0_st0_arr[1][7] <= 64'd16999845100481770868;
            ROM0_st0_arr[1][8] <= 64'd9335244255991628073;
            ROM0_st0_arr[1][9] <= 64'd12211248118271890408;
            ROM0_st0_arr[1][10] <= 64'd2714228989833617017;
            ROM0_st0_arr[1][11] <= 64'd2402649857173391264;
            ROM0_st0_arr[1][12] <= 64'd293230232171053580;
            ROM0_st0_arr[1][13] <= 64'd14925536787043292777;
            ROM0_st0_arr[1][14] <= 64'd1360553317005316379;
            ROM0_st0_arr[1][15] <= 64'd12653636911219766350;
            ROM0_st0_arr[2][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[2][1] <= 64'd3316608401227214173;
            ROM0_st0_arr[2][2] <= 64'd1191365957280576527;
            ROM0_st0_arr[2][3] <= 64'd2350022985419024820;
            ROM0_st0_arr[2][4] <= 64'd892617952471018716;
            ROM0_st0_arr[2][5] <= 64'd291466984857653829;
            ROM0_st0_arr[2][6] <= 64'd9195907541600953908;
            ROM0_st0_arr[2][7] <= 64'd13965188713800269600;
            ROM0_st0_arr[2][8] <= 64'd11671582227968848892;
            ROM0_st0_arr[2][9] <= 64'd5315256861805614728;
            ROM0_st0_arr[2][10] <= 64'd12995973883950975298;
            ROM0_st0_arr[2][11] <= 64'd2656329785076651114;
            ROM0_st0_arr[2][12] <= 64'd18166762397147179996;
            ROM0_st0_arr[2][13] <= 64'd18164872913915589634;
            ROM0_st0_arr[2][14] <= 64'd13678337806070825902;
            ROM0_st0_arr[2][15] <= 64'd558520734427554446;
            ROM0_st0_arr[3][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[3][1] <= 64'd15941224634913062555;
            ROM0_st0_arr[3][2] <= 64'd6226102851069492885;
            ROM0_st0_arr[3][3] <= 64'd6292042468883387737;
            ROM0_st0_arr[3][4] <= 64'd16466582063388455247;
            ROM0_st0_arr[3][5] <= 64'd8225018769583795339;
            ROM0_st0_arr[3][6] <= 64'd4512091954224483758;
            ROM0_st0_arr[3][7] <= 64'd8645835248368287205;
            ROM0_st0_arr[3][8] <= 64'd17111454092764159537;
            ROM0_st0_arr[3][9] <= 64'd2108312828726247716;
            ROM0_st0_arr[3][10] <= 64'd13801561118745443899;
            ROM0_st0_arr[3][11] <= 64'd12733692426302762269;
            ROM0_st0_arr[3][12] <= 64'd9260244138063238019;
            ROM0_st0_arr[3][13] <= 64'd13571746033574183535;
            ROM0_st0_arr[3][14] <= 64'd13490616479281253697;
            ROM0_st0_arr[3][15] <= 64'd8972334800401024692;
            ROM0_st0_arr[4][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[4][1] <= 64'd16450014459459345480;
            ROM0_st0_arr[4][2] <= 64'd9881659706905143497;
            ROM0_st0_arr[4][3] <= 64'd13975895267777782095;
            ROM0_st0_arr[4][4] <= 64'd8056503374861520973;
            ROM0_st0_arr[4][5] <= 64'd552255897587383266;
            ROM0_st0_arr[4][6] <= 64'd17714432001231460403;
            ROM0_st0_arr[4][7] <= 64'd8560833999250493496;
            ROM0_st0_arr[4][8] <= 64'd13855921957946101128;
            ROM0_st0_arr[4][9] <= 64'd1474323045092093876;
            ROM0_st0_arr[4][10] <= 64'd505394147197848886;
            ROM0_st0_arr[4][11] <= 64'd3136702942479751725;
            ROM0_st0_arr[4][12] <= 64'd7707559984774479304;
            ROM0_st0_arr[4][13] <= 64'd323638514611028602;
            ROM0_st0_arr[4][14] <= 64'd16000225301630982591;
            ROM0_st0_arr[4][15] <= 64'd3926266150091745462;
            ROM0_st0_arr[5][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[5][1] <= 64'd15982007350048747564;
            ROM0_st0_arr[5][2] <= 64'd6468410005745708178;
            ROM0_st0_arr[5][3] <= 64'd1047800296056156975;
            ROM0_st0_arr[5][4] <= 64'd4066165296528598587;
            ROM0_st0_arr[5][5] <= 64'd7997919790049200182;
            ROM0_st0_arr[5][6] <= 64'd17835182547887578391;
            ROM0_st0_arr[5][7] <= 64'd10559137563776343209;
            ROM0_st0_arr[5][8] <= 64'd2089344228083915210;
            ROM0_st0_arr[5][9] <= 64'd3385412779512615198;
            ROM0_st0_arr[5][10] <= 64'd16746206278156419730;
            ROM0_st0_arr[5][11] <= 64'd673168403760943276;
            ROM0_st0_arr[5][12] <= 64'd14186514604118539351;
            ROM0_st0_arr[5][13] <= 64'd4922790228527992930;
            ROM0_st0_arr[5][14] <= 64'd5251625098839442018;
            ROM0_st0_arr[5][15] <= 64'd9451369126729375126;
            ROM0_st0_arr[6][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[6][1] <= 64'd892902153545801848;
            ROM0_st0_arr[6][2] <= 64'd4304840548186534192;
            ROM0_st0_arr[6][3] <= 64'd13677550649392937527;
            ROM0_st0_arr[6][4] <= 64'd3621112023867626175;
            ROM0_st0_arr[6][5] <= 64'd7528509930910318757;
            ROM0_st0_arr[6][6] <= 64'd8758621768662845155;
            ROM0_st0_arr[6][7] <= 64'd15138477949936628362;
            ROM0_st0_arr[6][8] <= 64'd2849657757282217625;
            ROM0_st0_arr[6][9] <= 64'd13732447940012066702;
            ROM0_st0_arr[6][10] <= 64'd4367124966835549543;
            ROM0_st0_arr[6][11] <= 64'd7570866175719707247;
            ROM0_st0_arr[6][12] <= 64'd16100902212046155681;
            ROM0_st0_arr[6][13] <= 64'd3255920939831394824;
            ROM0_st0_arr[6][14] <= 64'd15879737847372079554;
            ROM0_st0_arr[6][15] <= 64'd13978578193994148753;
            ROM0_st0_arr[7][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[7][1] <= 64'd12915879621690710083;
            ROM0_st0_arr[7][2] <= 64'd5955555040728699654;
            ROM0_st0_arr[7][3] <= 64'd11199236800359540003;
            ROM0_st0_arr[7][4] <= 64'd16942058356233310568;
            ROM0_st0_arr[7][5] <= 64'd4915431680932952579;
            ROM0_st0_arr[7][6] <= 64'd12928550677510489252;
            ROM0_st0_arr[7][7] <= 64'd3302201367451394411;
            ROM0_st0_arr[7][8] <= 64'd7161233499657537350;
            ROM0_st0_arr[7][9] <= 64'd7719623134377957305;
            ROM0_st0_arr[7][10] <= 64'd15179656220160232506;
            ROM0_st0_arr[7][11] <= 64'd7717425068983310428;
            ROM0_st0_arr[7][12] <= 64'd2239853378139234600;
            ROM0_st0_arr[7][13] <= 64'd12758199090098265224;
            ROM0_st0_arr[7][14] <= 64'd6758255710041476138;
            ROM0_st0_arr[7][15] <= 64'd2008297874450139748;
            ROM0_st0_arr[8][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[8][1] <= 64'd16836943338755067060;
            ROM0_st0_arr[8][2] <= 64'd2439672451841033053;
            ROM0_st0_arr[8][3] <= 64'd811209873465104844;
            ROM0_st0_arr[8][4] <= 64'd18101933817957049782;
            ROM0_st0_arr[8][5] <= 64'd4680079369449503840;
            ROM0_st0_arr[8][6] <= 64'd11965081838267927603;
            ROM0_st0_arr[8][7] <= 64'd12265063152553980298;
            ROM0_st0_arr[8][8] <= 64'd1617487983075468259;
            ROM0_st0_arr[8][9] <= 64'd2302442326963614021;
            ROM0_st0_arr[8][10] <= 64'd6712673344879703542;
            ROM0_st0_arr[8][11] <= 64'd1775935601559311812;
            ROM0_st0_arr[8][12] <= 64'd18151767242567017453;
            ROM0_st0_arr[8][13] <= 64'd18128966925529969656;
            ROM0_st0_arr[8][14] <= 64'd8693490608450502988;
            ROM0_st0_arr[8][15] <= 64'd5483358938095204946;
            ROM0_st0_arr[9][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[9][1] <= 64'd4460188892089261596;
            ROM0_st0_arr[9][2] <= 64'd5087077863183075150;
            ROM0_st0_arr[9][3] <= 64'd13673491222243862709;
            ROM0_st0_arr[9][4] <= 64'd11264495381567969723;
            ROM0_st0_arr[9][5] <= 64'd1577020478793669798;
            ROM0_st0_arr[9][6] <= 64'd8594418532315835451;
            ROM0_st0_arr[9][7] <= 64'd11542928553390918846;
            ROM0_st0_arr[9][8] <= 64'd10062789913225546609;
            ROM0_st0_arr[9][9] <= 64'd16110920432432586900;
            ROM0_st0_arr[9][10] <= 64'd267975466523954734;
            ROM0_st0_arr[9][11] <= 64'd3923652581253579948;
            ROM0_st0_arr[9][12] <= 64'd12126496399462502852;
            ROM0_st0_arr[9][13] <= 64'd11711403565948912504;
            ROM0_st0_arr[9][14] <= 64'd16537066578843160879;
            ROM0_st0_arr[9][15] <= 64'd16622767333237920597;
            ROM0_st0_arr[10][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[10][1] <= 64'd8306858900184308299;
            ROM0_st0_arr[10][2] <= 64'd13767794918495523644;
            ROM0_st0_arr[10][3] <= 64'd15739227304438918407;
            ROM0_st0_arr[10][4] <= 64'd15281597592662976618;
            ROM0_st0_arr[10][5] <= 64'd13891151922390022198;
            ROM0_st0_arr[10][6] <= 64'd13959084736526763319;
            ROM0_st0_arr[10][7] <= 64'd1242666940968777068;
            ROM0_st0_arr[10][8] <= 64'd13966057335751391955;
            ROM0_st0_arr[10][9] <= 64'd10714610275495456146;
            ROM0_st0_arr[10][10] <= 64'd14403590891831793233;
            ROM0_st0_arr[10][11] <= 64'd8118143573377463433;
            ROM0_st0_arr[10][12] <= 64'd15635091652953775439;
            ROM0_st0_arr[10][13] <= 64'd6824554946361560998;
            ROM0_st0_arr[10][14] <= 64'd14736829215404272606;
            ROM0_st0_arr[10][15] <= 64'd17298582933948900223;
            ROM0_st0_arr[11][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[11][1] <= 64'd7533138519363761158;
            ROM0_st0_arr[11][2] <= 64'd1636326708996231348;
            ROM0_st0_arr[11][3] <= 64'd15372520741003543715;
            ROM0_st0_arr[11][4] <= 64'd16829584448654570394;
            ROM0_st0_arr[11][5] <= 64'd13824276422359892444;
            ROM0_st0_arr[11][6] <= 64'd9306920784263974807;
            ROM0_st0_arr[11][7] <= 64'd14966414557708197430;
            ROM0_st0_arr[11][8] <= 64'd5258157499736339221;
            ROM0_st0_arr[11][9] <= 64'd10012051443840883661;
            ROM0_st0_arr[11][10] <= 64'd13604302330065316728;
            ROM0_st0_arr[11][11] <= 64'd1829787159420351885;
            ROM0_st0_arr[11][12] <= 64'd319990789532844799;
            ROM0_st0_arr[11][13] <= 64'd2050533557548945054;
            ROM0_st0_arr[11][14] <= 64'd8880132830079482804;
            ROM0_st0_arr[11][15] <= 64'd2380361073813466337;
            ROM0_st0_arr[12][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[12][1] <= 64'd2048811532747770767;
            ROM0_st0_arr[12][2] <= 64'd8320561024393467379;
            ROM0_st0_arr[12][3] <= 64'd5211666985007417987;
            ROM0_st0_arr[12][4] <= 64'd11866900833167961951;
            ROM0_st0_arr[12][5] <= 64'd7151135148549474616;
            ROM0_st0_arr[12][6] <= 64'd219715944850706020;
            ROM0_st0_arr[12][7] <= 64'd6381770425018462736;
            ROM0_st0_arr[12][8] <= 64'd5970679186843280180;
            ROM0_st0_arr[12][9] <= 64'd7143498643723256195;
            ROM0_st0_arr[12][10] <= 64'd1956488404144772298;
            ROM0_st0_arr[12][11] <= 64'd5619747107484077139;
            ROM0_st0_arr[12][12] <= 64'd527917044300707521;
            ROM0_st0_arr[12][13] <= 64'd3318798955808550409;
            ROM0_st0_arr[12][14] <= 64'd4358843149513399777;
            ROM0_st0_arr[12][15] <= 64'd11473360703482113395;
            ROM0_st0_arr[13][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[13][1] <= 64'd12432417682878015040;
            ROM0_st0_arr[13][2] <= 64'd3955739673572204771;
            ROM0_st0_arr[13][3] <= 64'd8992488188073208194;
            ROM0_st0_arr[13][4] <= 64'd7231027521189447218;
            ROM0_st0_arr[13][5] <= 64'd8055849936219707510;
            ROM0_st0_arr[13][6] <= 64'd796752505033298578;
            ROM0_st0_arr[13][7] <= 64'd1520483667984614851;
            ROM0_st0_arr[13][8] <= 64'd14894687694104923508;
            ROM0_st0_arr[13][9] <= 64'd11015921181254749521;
            ROM0_st0_arr[13][10] <= 64'd7689958724620230199;
            ROM0_st0_arr[13][11] <= 64'd3558381302344981306;
            ROM0_st0_arr[13][12] <= 64'd2359814614780534944;
            ROM0_st0_arr[13][13] <= 64'd1046803206103297723;
            ROM0_st0_arr[13][14] <= 64'd16693924160465396879;
            ROM0_st0_arr[13][15] <= 64'd14591813889413309792;
            ROM0_st0_arr[14][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[14][1] <= 64'd16126949464588608127;
            ROM0_st0_arr[14][2] <= 64'd17078700769474680244;
            ROM0_st0_arr[14][3] <= 64'd12577868261904608354;
            ROM0_st0_arr[14][4] <= 64'd8749721333104439875;
            ROM0_st0_arr[14][5] <= 64'd16115008190553353689;
            ROM0_st0_arr[14][6] <= 64'd5858496545464991344;
            ROM0_st0_arr[14][7] <= 64'd126526973274617528;
            ROM0_st0_arr[14][8] <= 64'd14755250061178960331;
            ROM0_st0_arr[14][9] <= 64'd2950081247540242882;
            ROM0_st0_arr[14][10] <= 64'd1638845449206124627;
            ROM0_st0_arr[14][11] <= 64'd5167612594998720597;
            ROM0_st0_arr[14][12] <= 64'd13668493220787483110;
            ROM0_st0_arr[14][13] <= 64'd7737503417762794307;
            ROM0_st0_arr[14][14] <= 64'd18260109989201046983;
            ROM0_st0_arr[14][15] <= 64'd9185289083725472784;
            ROM0_st0_arr[15][0] <= 64'd17293822565076172801;
            ROM0_st0_arr[15][1] <= 64'd662880509164891295;
            ROM0_st0_arr[15][2] <= 64'd14962411951571283646;
            ROM0_st0_arr[15][3] <= 64'd7586481955073758662;
            ROM0_st0_arr[15][4] <= 64'd14298533999211558888;
            ROM0_st0_arr[15][5] <= 64'd7986826120987974572;
            ROM0_st0_arr[15][6] <= 64'd4892492172216047440;
            ROM0_st0_arr[15][7] <= 64'd303693874776087318;
            ROM0_st0_arr[15][8] <= 64'd2939983354724710425;
            ROM0_st0_arr[15][9] <= 64'd8633471479223067074;
            ROM0_st0_arr[15][10] <= 64'd16302940337222946449;
            ROM0_st0_arr[15][11] <= 64'd11899329780723059891;
            ROM0_st0_arr[15][12] <= 64'd4046475262271886735;
            ROM0_st0_arr[15][13] <= 64'd16855513577843145672;
            ROM0_st0_arr[15][14] <= 64'd6747459861404804573;
            ROM0_st0_arr[15][15] <= 64'd17850599548321437946;

            ROM0_st1_arr[0][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[0][1] <= 64'd10405021248184179819;
            ROM0_st1_arr[0][2] <= 64'd18357364935460720835;
            ROM0_st1_arr[0][3] <= 64'd7524045725815612048;
            ROM0_st1_arr[0][4] <= 64'd14020921120480921444;
            ROM0_st1_arr[0][5] <= 64'd4567431763498152711;
            ROM0_st1_arr[0][6] <= 64'd16649986813178928548;
            ROM0_st1_arr[0][7] <= 64'd6260718610716965298;
            ROM0_st1_arr[0][8] <= 64'd14265650877534657191;
            ROM0_st1_arr[0][9] <= 64'd2205622138389660681;
            ROM0_st1_arr[0][10] <= 64'd11557582455713433260;
            ROM0_st1_arr[0][11] <= 64'd1274458201404381182;
            ROM0_st1_arr[0][12] <= 64'd8995418809887038361;
            ROM0_st1_arr[0][13] <= 64'd13028762822951290503;
            ROM0_st1_arr[0][14] <= 64'd5332075283400248574;
            ROM0_st1_arr[0][15] <= 64'd15461929222870183236;
            ROM0_st1_arr[1][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[1][1] <= 64'd6427090851680715034;
            ROM0_st1_arr[1][2] <= 64'd7019646305631508202;
            ROM0_st1_arr[1][3] <= 64'd3543018840566806211;
            ROM0_st1_arr[1][4] <= 64'd13482549406713562221;
            ROM0_st1_arr[1][5] <= 64'd6636031775788163037;
            ROM0_st1_arr[1][6] <= 64'd6686419642167453063;
            ROM0_st1_arr[1][7] <= 64'd14975756600363089480;
            ROM0_st1_arr[1][8] <= 64'd11018083872338033302;
            ROM0_st1_arr[1][9] <= 64'd12397375900707528775;
            ROM0_st1_arr[1][10] <= 64'd3499557463425346777;
            ROM0_st1_arr[1][11] <= 64'd14664756014577757064;
            ROM0_st1_arr[1][12] <= 64'd18257403526048309240;
            ROM0_st1_arr[1][13] <= 64'd772415948059296082;
            ROM0_st1_arr[1][14] <= 64'd5302101404170755547;
            ROM0_st1_arr[1][15] <= 64'd3562911137331613973;
            ROM0_st1_arr[2][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[2][1] <= 64'd2243039484195993191;
            ROM0_st1_arr[2][2] <= 64'd8132681561913633117;
            ROM0_st1_arr[2][3] <= 64'd2021821058377181664;
            ROM0_st1_arr[2][4] <= 64'd10157216646538189283;
            ROM0_st1_arr[2][5] <= 64'd9171185784906045668;
            ROM0_st1_arr[2][6] <= 64'd4305380472265991609;
            ROM0_st1_arr[2][7] <= 64'd2211928315324603342;
            ROM0_st1_arr[2][8] <= 64'd6168910713355981590;
            ROM0_st1_arr[2][9] <= 64'd17878253867428005688;
            ROM0_st1_arr[2][10] <= 64'd13760077253876019195;
            ROM0_st1_arr[2][11] <= 64'd52960884282847133;
            ROM0_st1_arr[2][12] <= 64'd14332178914760844213;
            ROM0_st1_arr[2][13] <= 64'd1138901487548130847;
            ROM0_st1_arr[2][14] <= 64'd4303843542009117362;
            ROM0_st1_arr[2][15] <= 64'd14035891226182752717;
            ROM0_st1_arr[3][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[3][1] <= 64'd15985486925786043797;
            ROM0_st1_arr[3][2] <= 64'd17023943044813816274;
            ROM0_st1_arr[3][3] <= 64'd8274139857233974205;
            ROM0_st1_arr[3][4] <= 64'd12759702089327230191;
            ROM0_st1_arr[3][5] <= 64'd13103308231302819623;
            ROM0_st1_arr[3][6] <= 64'd5734663407885852338;
            ROM0_st1_arr[3][7] <= 64'd5852366706506290297;
            ROM0_st1_arr[3][8] <= 64'd6244679043965076148;
            ROM0_st1_arr[3][9] <= 64'd9348487763318866904;
            ROM0_st1_arr[3][10] <= 64'd14858417106656830991;
            ROM0_st1_arr[3][11] <= 64'd7988408224489878966;
            ROM0_st1_arr[3][12] <= 64'd13257964703471134012;
            ROM0_st1_arr[3][13] <= 64'd6177496660492614933;
            ROM0_st1_arr[3][14] <= 64'd16752761998819501770;
            ROM0_st1_arr[3][15] <= 64'd9706686830946461896;
            ROM0_st1_arr[4][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[4][1] <= 64'd15961793146812735399;
            ROM0_st1_arr[4][2] <= 64'd577857301137234877;
            ROM0_st1_arr[4][3] <= 64'd5047087551566044369;
            ROM0_st1_arr[4][4] <= 64'd9929356652858941593;
            ROM0_st1_arr[4][5] <= 64'd3246800698745713157;
            ROM0_st1_arr[4][6] <= 64'd17827717081112796515;
            ROM0_st1_arr[4][7] <= 64'd13714931867796837460;
            ROM0_st1_arr[4][8] <= 64'd14890406446337395446;
            ROM0_st1_arr[4][9] <= 64'd3803362446657989762;
            ROM0_st1_arr[4][10] <= 64'd18183312823727473992;
            ROM0_st1_arr[4][11] <= 64'd1982229535856330968;
            ROM0_st1_arr[4][12] <= 64'd8713636547823424534;
            ROM0_st1_arr[4][13] <= 64'd11451956292395797655;
            ROM0_st1_arr[4][14] <= 64'd14812248543932043928;
            ROM0_st1_arr[4][15] <= 64'd5431774702940624359;
            ROM0_st1_arr[5][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[5][1] <= 64'd2577671089079286439;
            ROM0_st1_arr[5][2] <= 64'd11995993822027828645;
            ROM0_st1_arr[5][3] <= 64'd3042797204296855209;
            ROM0_st1_arr[5][4] <= 64'd13347457330830597389;
            ROM0_st1_arr[5][5] <= 64'd886530956755740804;
            ROM0_st1_arr[5][6] <= 64'd8746457548859571803;
            ROM0_st1_arr[5][7] <= 64'd13098305493279876251;
            ROM0_st1_arr[5][8] <= 64'd15331777707844533717;
            ROM0_st1_arr[5][9] <= 64'd8532094430781013622;
            ROM0_st1_arr[5][10] <= 64'd15718604359612274874;
            ROM0_st1_arr[5][11] <= 64'd2957922565978088898;
            ROM0_st1_arr[5][12] <= 64'd1823625798562030396;
            ROM0_st1_arr[5][13] <= 64'd8095339948653323243;
            ROM0_st1_arr[5][14] <= 64'd13792745165838085667;
            ROM0_st1_arr[5][15] <= 64'd8390199040176256858;
            ROM0_st1_arr[6][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[6][1] <= 64'd14618045663912337671;
            ROM0_st1_arr[6][2] <= 64'd8231607757048583003;
            ROM0_st1_arr[6][3] <= 64'd18127352228187063615;
            ROM0_st1_arr[6][4] <= 64'd7050613204414151038;
            ROM0_st1_arr[6][5] <= 64'd13505419564446567997;
            ROM0_st1_arr[6][6] <= 64'd6444142060334423532;
            ROM0_st1_arr[6][7] <= 64'd6056783327295541961;
            ROM0_st1_arr[6][8] <= 64'd5813278871091589641;
            ROM0_st1_arr[6][9] <= 64'd2705129707231313014;
            ROM0_st1_arr[6][10] <= 64'd18219804770780039846;
            ROM0_st1_arr[6][11] <= 64'd17018430414050656351;
            ROM0_st1_arr[6][12] <= 64'd1514724346930200648;
            ROM0_st1_arr[6][13] <= 64'd11268495472790879713;
            ROM0_st1_arr[6][14] <= 64'd7351163212087983469;
            ROM0_st1_arr[6][15] <= 64'd16840078676440068511;
            ROM0_st1_arr[7][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[7][1] <= 64'd1596492687493210785;
            ROM0_st1_arr[7][2] <= 64'd4922147659447635961;
            ROM0_st1_arr[7][3] <= 64'd7756028884659941004;
            ROM0_st1_arr[7][4] <= 64'd3538440868305609356;
            ROM0_st1_arr[7][5] <= 64'd7364503734003393836;
            ROM0_st1_arr[7][6] <= 64'd16693836776352278179;
            ROM0_st1_arr[7][7] <= 64'd16433977088157531717;
            ROM0_st1_arr[7][8] <= 64'd2503240902400619832;
            ROM0_st1_arr[7][9] <= 64'd212845868149098608;
            ROM0_st1_arr[7][10] <= 64'd8897028431426394426;
            ROM0_st1_arr[7][11] <= 64'd13584388978012141423;
            ROM0_st1_arr[7][12] <= 64'd14469777167815336543;
            ROM0_st1_arr[7][13] <= 64'd8485054302324926805;
            ROM0_st1_arr[7][14] <= 64'd14144279383711108454;
            ROM0_st1_arr[7][15] <= 64'd14580225699501226437;
            ROM0_st1_arr[8][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[8][1] <= 64'd12231327714635046031;
            ROM0_st1_arr[8][2] <= 64'd17573023920830506386;
            ROM0_st1_arr[8][3] <= 64'd5234279963735994814;
            ROM0_st1_arr[8][4] <= 64'd17760117485926407451;
            ROM0_st1_arr[8][5] <= 64'd6670618412913399791;
            ROM0_st1_arr[8][6] <= 64'd1682237559320119303;
            ROM0_st1_arr[8][7] <= 64'd466014321377454543;
            ROM0_st1_arr[8][8] <= 64'd16101787921637751596;
            ROM0_st1_arr[8][9] <= 64'd4600071385601631992;
            ROM0_st1_arr[8][10] <= 64'd599846385479352366;
            ROM0_st1_arr[8][11] <= 64'd15735181537912819138;
            ROM0_st1_arr[8][12] <= 64'd4616746788718433830;
            ROM0_st1_arr[8][13] <= 64'd15783751702225169603;
            ROM0_st1_arr[8][14] <= 64'd764617379449676960;
            ROM0_st1_arr[8][15] <= 64'd11886034584718758091;
            ROM0_st1_arr[9][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[9][1] <= 64'd7393566483642163708;
            ROM0_st1_arr[9][2] <= 64'd10477086511661121738;
            ROM0_st1_arr[9][3] <= 64'd986485908852701152;
            ROM0_st1_arr[9][4] <= 64'd3403476374447959414;
            ROM0_st1_arr[9][5] <= 64'd12122422949187998102;
            ROM0_st1_arr[9][6] <= 64'd13805399445681343821;
            ROM0_st1_arr[9][7] <= 64'd7214158157271938108;
            ROM0_st1_arr[9][8] <= 64'd12430546111446936852;
            ROM0_st1_arr[9][9] <= 64'd15406786089292215038;
            ROM0_st1_arr[9][10] <= 64'd10259871632647442319;
            ROM0_st1_arr[9][11] <= 64'd12433442803623597191;
            ROM0_st1_arr[9][12] <= 64'd4077883895070941012;
            ROM0_st1_arr[9][13] <= 64'd12743382161634612512;
            ROM0_st1_arr[9][14] <= 64'd12857162286965609626;
            ROM0_st1_arr[9][15] <= 64'd6665383956248282420;
            ROM0_st1_arr[10][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[10][1] <= 64'd11205937175358949927;
            ROM0_st1_arr[10][2] <= 64'd7653601283080393651;
            ROM0_st1_arr[10][3] <= 64'd8824795755142539266;
            ROM0_st1_arr[10][4] <= 64'd7504718318566677644;
            ROM0_st1_arr[10][5] <= 64'd8772840058683537643;
            ROM0_st1_arr[10][6] <= 64'd14374058049885246184;
            ROM0_st1_arr[10][7] <= 64'd4095992279035047971;
            ROM0_st1_arr[10][8] <= 64'd5570380238700699212;
            ROM0_st1_arr[10][9] <= 64'd11844904009531608751;
            ROM0_st1_arr[10][10] <= 64'd2107449965496882632;
            ROM0_st1_arr[10][11] <= 64'd3592154860391298583;
            ROM0_st1_arr[10][12] <= 64'd3857737680918341153;
            ROM0_st1_arr[10][13] <= 64'd14085532411580104904;
            ROM0_st1_arr[10][14] <= 64'd6544182290997896124;
            ROM0_st1_arr[10][15] <= 64'd12853323143796126480;
            ROM0_st1_arr[11][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[11][1] <= 64'd5803064664561253546;
            ROM0_st1_arr[11][2] <= 64'd16352222879643494849;
            ROM0_st1_arr[11][3] <= 64'd4967227718261905131;
            ROM0_st1_arr[11][4] <= 64'd15511260990217806155;
            ROM0_st1_arr[11][5] <= 64'd17656006751039262143;
            ROM0_st1_arr[11][6] <= 64'd1848875070904128459;
            ROM0_st1_arr[11][7] <= 64'd4542768994119092665;
            ROM0_st1_arr[11][8] <= 64'd3371727321785536135;
            ROM0_st1_arr[11][9] <= 64'd14271832993747149179;
            ROM0_st1_arr[11][10] <= 64'd3378373609003891255;
            ROM0_st1_arr[11][11] <= 64'd5123107541484101187;
            ROM0_st1_arr[11][12] <= 64'd6328949293972979137;
            ROM0_st1_arr[11][13] <= 64'd9362946477935208725;
            ROM0_st1_arr[11][14] <= 64'd2574791057574424200;
            ROM0_st1_arr[11][15] <= 64'd12485402889892278751;
            ROM0_st1_arr[12][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[12][1] <= 64'd10991581649380563330;
            ROM0_st1_arr[12][2] <= 64'd4913568270759875178;
            ROM0_st1_arr[12][3] <= 64'd17812913537642853032;
            ROM0_st1_arr[12][4] <= 64'd3341503289287630222;
            ROM0_st1_arr[12][5] <= 64'd354034030843946954;
            ROM0_st1_arr[12][6] <= 64'd2450444360701235770;
            ROM0_st1_arr[12][7] <= 64'd10132164321287060717;
            ROM0_st1_arr[12][8] <= 64'd1964929393189321158;
            ROM0_st1_arr[12][9] <= 64'd10500707696816686377;
            ROM0_st1_arr[12][10] <= 64'd1815514389076355800;
            ROM0_st1_arr[12][11] <= 64'd12961593949203426608;
            ROM0_st1_arr[12][12] <= 64'd13368991143379397903;
            ROM0_st1_arr[12][13] <= 64'd1606969135698904138;
            ROM0_st1_arr[12][14] <= 64'd371208358915902681;
            ROM0_st1_arr[12][15] <= 64'd15592187738737441198;
            ROM0_st1_arr[13][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[13][1] <= 64'd11200708556532648470;
            ROM0_st1_arr[13][2] <= 64'd2718599284101323773;
            ROM0_st1_arr[13][3] <= 64'd11216836580702018198;
            ROM0_st1_arr[13][4] <= 64'd2928170683958478459;
            ROM0_st1_arr[13][5] <= 64'd2251978001938448667;
            ROM0_st1_arr[13][6] <= 64'd9462924945156934259;
            ROM0_st1_arr[13][7] <= 64'd248155003269738165;
            ROM0_st1_arr[13][8] <= 64'd1698680234739034137;
            ROM0_st1_arr[13][9] <= 64'd14579436371013092868;
            ROM0_st1_arr[13][10] <= 64'd2610748826247181876;
            ROM0_st1_arr[13][11] <= 64'd14182472021891143239;
            ROM0_st1_arr[13][12] <= 64'd18406257898496282323;
            ROM0_st1_arr[13][13] <= 64'd12911010253573340831;
            ROM0_st1_arr[13][14] <= 64'd7292885344072883191;
            ROM0_st1_arr[13][15] <= 64'd2017160558257493603;
            ROM0_st1_arr[14][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[14][1] <= 64'd1789205669093589884;
            ROM0_st1_arr[14][2] <= 64'd14580161660266615730;
            ROM0_st1_arr[14][3] <= 64'd8164886603416501794;
            ROM0_st1_arr[14][4] <= 64'd3983014276289321098;
            ROM0_st1_arr[14][5] <= 64'd417489998409971940;
            ROM0_st1_arr[14][6] <= 64'd4952215906414302448;
            ROM0_st1_arr[14][7] <= 64'd14439733804589825819;
            ROM0_st1_arr[14][8] <= 64'd7179217523447274592;
            ROM0_st1_arr[14][9] <= 64'd12548826928377459663;
            ROM0_st1_arr[14][10] <= 64'd13647972985579765393;
            ROM0_st1_arr[14][11] <= 64'd943441632390584557;
            ROM0_st1_arr[14][12] <= 64'd4270416978261640546;
            ROM0_st1_arr[14][13] <= 64'd17562407657325825658;
            ROM0_st1_arr[14][14] <= 64'd13168548641635907169;
            ROM0_st1_arr[14][15] <= 64'd7853879266118494086;
            ROM0_st1_arr[15][0] <= 64'd17293822565076172801;
            ROM0_st1_arr[15][1] <= 64'd9486657212549813622;
            ROM0_st1_arr[15][2] <= 64'd32726893590173273;
            ROM0_st1_arr[15][3] <= 64'd14673542420584572300;
            ROM0_st1_arr[15][4] <= 64'd16959839522054718695;
            ROM0_st1_arr[15][5] <= 64'd5853998566064948942;
            ROM0_st1_arr[15][6] <= 64'd3815315886781762860;
            ROM0_st1_arr[15][7] <= 64'd6273129929571326275;
            ROM0_st1_arr[15][8] <= 64'd9111196760903428495;
            ROM0_st1_arr[15][9] <= 64'd10365740339457113609;
            ROM0_st1_arr[15][10] <= 64'd10154747285893383053;
            ROM0_st1_arr[15][11] <= 64'd9829856391104209805;
            ROM0_st1_arr[15][12] <= 64'd6031586691482439418;
            ROM0_st1_arr[15][13] <= 64'd16121882724449528061;
            ROM0_st1_arr[15][14] <= 64'd6254766350509124677;
            ROM0_st1_arr[15][15] <= 64'd10797241297349275918;

            ROM0_st2_arr[0][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[0][1] <= 64'd12154600967831981241;
            ROM0_st2_arr[0][2] <= 64'd14276274543166211387;
            ROM0_st2_arr[0][3] <= 64'd418881448437566951;
            ROM0_st2_arr[0][4] <= 64'd18158518091376492545;
            ROM0_st2_arr[0][5] <= 64'd118607460926999667;
            ROM0_st2_arr[0][6] <= 64'd4889317495851452527;
            ROM0_st2_arr[0][7] <= 64'd2272940007883440574;
            ROM0_st2_arr[0][8] <= 64'd2199023255552;
            ROM0_st2_arr[0][9] <= 64'd10069193652868617379;
            ROM0_st2_arr[0][10] <= 64'd16801025490767711121;
            ROM0_st2_arr[0][11] <= 64'd17225010883624785699;
            ROM0_st2_arr[0][12] <= 64'd36029346766389248;
            ROM0_st2_arr[0][13] <= 64'd2713927885141610691;
            ROM0_st2_arr[0][14] <= 64'd14706877084432893115;
            ROM0_st2_arr[0][15] <= 64'd12940073958180608858;
            ROM0_st2_arr[1][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[1][1] <= 64'd418881448437566951;
            ROM0_st2_arr[1][2] <= 64'd4889317495851452527;
            ROM0_st2_arr[1][3] <= 64'd10069193652868617379;
            ROM0_st2_arr[1][4] <= 64'd36029346766389248;
            ROM0_st2_arr[1][5] <= 64'd12940073958180608858;
            ROM0_st2_arr[1][6] <= 64'd16782525399254597868;
            ROM0_st2_arr[1][7] <= 64'd14697895938737762511;
            ROM0_st2_arr[1][8] <= 64'd18446744035054845953;
            ROM0_st2_arr[1][9] <= 64'd9818922367904463524;
            ROM0_st2_arr[1][10] <= 64'd16775797234547305966;
            ROM0_st2_arr[1][11] <= 64'd3781487518361002985;
            ROM0_st2_arr[1][12] <= 64'd18446673701744164865;
            ROM0_st2_arr[1][13] <= 64'd16438693553069120169;
            ROM0_st2_arr[1][14] <= 64'd5115687388739336161;
            ROM0_st2_arr[1][15] <= 64'd17569204722331893322;
            ROM0_st2_arr[2][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[2][1] <= 64'd118607460926999667;
            ROM0_st2_arr[2][2] <= 64'd16801025490767711121;
            ROM0_st2_arr[2][3] <= 64'd12940073958180608858;
            ROM0_st2_arr[2][4] <= 64'd4503530906845184;
            ROM0_st2_arr[2][5] <= 64'd9930732012135028654;
            ROM0_st2_arr[2][6] <= 64'd16775797234547305966;
            ROM0_st2_arr[2][7] <= 64'd2418535265313493493;
            ROM0_st2_arr[2][8] <= 64'd536870912;
            ROM0_st2_arr[2][9] <= 64'd17569204722331893322;
            ROM0_st2_arr[2][10] <= 64'd17387991853842663593;
            ROM0_st2_arr[2][11] <= 64'd11560590832702013078;
            ROM0_st2_arr[2][12] <= 64'd18446743931973533729;
            ROM0_st2_arr[2][13] <= 64'd13939564058192504755;
            ROM0_st2_arr[2][14] <= 64'd12391532617460140695;
            ROM0_st2_arr[2][15] <= 64'd5668024148486473211;
            ROM0_st2_arr[3][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[3][1] <= 64'd2272940007883440574;
            ROM0_st2_arr[3][2] <= 64'd14706877084432893115;
            ROM0_st2_arr[3][3] <= 64'd14697895938737762511;
            ROM0_st2_arr[3][4] <= 64'd18446181110871359489;
            ROM0_st2_arr[3][5] <= 64'd2418535265313493493;
            ROM0_st2_arr[3][6] <= 64'd5115687388739336161;
            ROM0_st2_arr[3][7] <= 64'd11758359676994327409;
            ROM0_st2_arr[3][8] <= 64'd18446744069406195713;
            ROM0_st2_arr[3][9] <= 64'd15480652140551887064;
            ROM0_st2_arr[3][10] <= 64'd12391532617460140695;
            ROM0_st2_arr[3][11] <= 64'd1976865992950664020;
            ROM0_st2_arr[3][12] <= 64'd1152921504606842880;
            ROM0_st2_arr[3][13] <= 64'd16917029311671468777;
            ROM0_st2_arr[3][14] <= 64'd7073470201911047317;
            ROM0_st2_arr[3][15] <= 64'd6602944137259479215;
            ROM0_st2_arr[4][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[4][1] <= 64'd10069193652868617379;
            ROM0_st2_arr[4][2] <= 64'd16782525399254597868;
            ROM0_st2_arr[4][3] <= 64'd9818922367904463524;
            ROM0_st2_arr[4][4] <= 64'd18446673701744164865;
            ROM0_st2_arr[4][5] <= 64'd17569204722331893322;
            ROM0_st2_arr[4][6] <= 64'd151907467378121323;
            ROM0_st2_arr[4][7] <= 64'd15480652140551887064;
            ROM0_st2_arr[4][8] <= 64'd131072;
            ROM0_st2_arr[4][9] <= 64'd14481943491905488994;
            ROM0_st2_arr[4][10] <= 64'd4465369883443651344;
            ROM0_st2_arr[4][11] <= 64'd4318401330473269126;
            ROM0_st2_arr[4][12] <= 64'd2251799813685256;
            ROM0_st2_arr[4][13] <= 64'd6025271986410849717;
            ROM0_st2_arr[4][14] <= 64'd16225692241432132747;
            ROM0_st2_arr[4][15] <= 64'd7159872751042635062;
            ROM0_st2_arr[5][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[5][1] <= 64'd17225010883624785699;
            ROM0_st2_arr[5][2] <= 64'd13470432090103656415;
            ROM0_st2_arr[5][3] <= 64'd3781487518361002985;
            ROM0_st2_arr[5][4] <= 64'd8796227237888;
            ROM0_st2_arr[5][5] <= 64'd11560590832702013078;
            ROM0_st2_arr[5][6] <= 64'd11545758046752426462;
            ROM0_st2_arr[5][7] <= 64'd1976865992950664020;
            ROM0_st2_arr[5][8] <= 64'd18446744069414582273;
            ROM0_st2_arr[5][9] <= 64'd4318401330473269126;
            ROM0_st2_arr[5][10] <= 64'd13020108504974810489;
            ROM0_st2_arr[5][11] <= 64'd13443656673831655998;
            ROM0_st2_arr[5][12] <= 64'd18158509295283470337;
            ROM0_st2_arr[5][13] <= 64'd4895803518339076152;
            ROM0_st2_arr[5][14] <= 64'd11321187709614116894;
            ROM0_st2_arr[5][15] <= 64'd7020314776661527992;
            ROM0_st2_arr[6][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[6][1] <= 64'd2713927885141610691;
            ROM0_st2_arr[6][2] <= 64'd4637400370145003474;
            ROM0_st2_arr[6][3] <= 64'd16438693553069120169;
            ROM0_st2_arr[6][4] <= 64'd1099494850304;
            ROM0_st2_arr[6][5] <= 64'd13939564058192504755;
            ROM0_st2_arr[6][6] <= 64'd827331699260490933;
            ROM0_st2_arr[6][7] <= 64'd16917029311671468777;
            ROM0_st2_arr[6][8] <= 64'd32;
            ROM0_st2_arr[6][9] <= 64'd6025271986410849717;
            ROM0_st2_arr[6][10] <= 64'd13165748629174985600;
            ROM0_st2_arr[6][11] <= 64'd4895803518339076152;
            ROM0_st2_arr[6][12] <= 64'd562941363355648;
            ROM0_st2_arr[6][13] <= 64'd16613587000532886654;
            ROM0_st2_arr[6][14] <= 64'd17765460494250502634;
            ROM0_st2_arr[6][15] <= 64'd9996039020351967275;
            ROM0_st2_arr[7][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[7][1] <= 64'd12940073958180608858;
            ROM0_st2_arr[7][2] <= 64'd16775797234547305966;
            ROM0_st2_arr[7][3] <= 64'd17569204722331893322;
            ROM0_st2_arr[7][4] <= 64'd18446743931973533729;
            ROM0_st2_arr[7][5] <= 64'd5668024148486473211;
            ROM0_st2_arr[7][6] <= 64'd4465369883443651344;
            ROM0_st2_arr[7][7] <= 64'd6602944137259479215;
            ROM0_st2_arr[7][8] <= 64'd9223372034707292160;
            ROM0_st2_arr[7][9] <= 64'd7159872751042635062;
            ROM0_st2_arr[7][10] <= 64'd13367574678938226840;
            ROM0_st2_arr[7][11] <= 64'd7020314776661527992;
            ROM0_st2_arr[7][12] <= 64'd1099528404736;
            ROM0_st2_arr[7][13] <= 64'd9996039020351967275;
            ROM0_st2_arr[7][14] <= 64'd1170529071279957890;
            ROM0_st2_arr[7][15] <= 64'd2516679110167919243;
            ROM0_st2_arr[8][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[8][1] <= 64'd16239215796699989454;
            ROM0_st2_arr[8][2] <= 64'd12419909588359173629;
            ROM0_st2_arr[8][3] <= 64'd15238420318963429305;
            ROM0_st2_arr[8][4] <= 64'd18446744052234977285;
            ROM0_st2_arr[8][5] <= 64'd16217235531541203655;
            ROM0_st2_arr[8][6] <= 64'd6240510758973793805;
            ROM0_st2_arr[8][7] <= 64'd2936745668635964057;
            ROM0_st2_arr[8][8] <= 64'd18302628881372282881;
            ROM0_st2_arr[8][9] <= 64'd6641587991941144762;
            ROM0_st2_arr[8][10] <= 64'd8470017724575365824;
            ROM0_st2_arr[8][11] <= 64'd18045703600608189944;
            ROM0_st2_arr[8][12] <= 64'd9223372032559841281;
            ROM0_st2_arr[8][13] <= 64'd4332997450119473497;
            ROM0_st2_arr[8][14] <= 64'd7697592870902193346;
            ROM0_st2_arr[8][15] <= 64'd16507994269317256788;
            ROM0_st2_arr[9][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[9][1] <= 64'd11234439644667675337;
            ROM0_st2_arr[9][2] <= 64'd8724666157214819649;
            ROM0_st2_arr[9][3] <= 64'd9595091699185839754;
            ROM0_st2_arr[9][4] <= 64'd9223372036854808576;
            ROM0_st2_arr[9][5] <= 64'd8254373971510759366;
            ROM0_st2_arr[9][6] <= 64'd5942314925871800366;
            ROM0_st2_arr[9][7] <= 64'd15182065057696283114;
            ROM0_st2_arr[9][8] <= 64'd2251799813160960;
            ROM0_st2_arr[9][9] <= 64'd7219845934194655807;
            ROM0_st2_arr[9][10] <= 64'd11548203476806380366;
            ROM0_st2_arr[9][11] <= 64'd4953233573984427337;
            ROM0_st2_arr[9][12] <= 64'd18428729670905102273;
            ROM0_st2_arr[9][13] <= 64'd16340952018638106489;
            ROM0_st2_arr[9][14] <= 64'd1645718578646873200;
            ROM0_st2_arr[9][15] <= 64'd17624458064366113348;
            ROM0_st2_arr[10][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[10][1] <= 64'd14697895938737762511;
            ROM0_st2_arr[10][2] <= 64'd5115687388739336161;
            ROM0_st2_arr[10][3] <= 64'd15480652140551887064;
            ROM0_st2_arr[10][4] <= 64'd1152921504606842880;
            ROM0_st2_arr[10][5] <= 64'd6602944137259479215;
            ROM0_st2_arr[10][6] <= 64'd16225692241432132747;
            ROM0_st2_arr[10][7] <= 64'd13682341403837213413;
            ROM0_st2_arr[10][8] <= 64'd18446708885042503681;
            ROM0_st2_arr[10][9] <= 64'd2189760912533326910;
            ROM0_st2_arr[10][10] <= 64'd1170529071279957890;
            ROM0_st2_arr[10][11] <= 64'd5643482763792491001;
            ROM0_st2_arr[10][12] <= 64'd2305878193048911872;
            ROM0_st2_arr[10][13] <= 64'd2207528272714594867;
            ROM0_st2_arr[10][14] <= 64'd9722077912199764672;
            ROM0_st2_arr[10][15] <= 64'd12265408184257183405;
            ROM0_st2_arr[11][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[11][1] <= 64'd17834768629622199802;
            ROM0_st2_arr[11][2] <= 64'd12996475468101930825;
            ROM0_st2_arr[11][3] <= 64'd13561337937994272377;
            ROM0_st2_arr[11][4] <= 64'd18302628881338727937;
            ROM0_st2_arr[11][5] <= 64'd1661907235718972450;
            ROM0_st2_arr[11][6] <= 64'd13313749361279891624;
            ROM0_st2_arr[11][7] <= 64'd5853027518870524662;
            ROM0_st2_arr[11][8] <= 64'd549755813760;
            ROM0_st2_arr[11][9] <= 64'd5381740272616182881;
            ROM0_st2_arr[11][10] <= 64'd6519596376689022014;
            ROM0_st2_arr[11][11] <= 64'd7670688024331825335;
            ROM0_st2_arr[11][12] <= 64'd18442240538507739137;
            ROM0_st2_arr[11][13] <= 64'd8223871192367387883;
            ROM0_st2_arr[11][14] <= 64'd6900986022662157859;
            ROM0_st2_arr[11][15] <= 64'd16760055257485814698;
            ROM0_st2_arr[12][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[12][1] <= 64'd9930732012135028654;
            ROM0_st2_arr[12][2] <= 64'd17387991853842663593;
            ROM0_st2_arr[12][3] <= 64'd5668024148486473211;
            ROM0_st2_arr[12][4] <= 64'd18428729670905102401;
            ROM0_st2_arr[12][5] <= 64'd17497884381998586985;
            ROM0_st2_arr[12][6] <= 64'd13367574678938226840;
            ROM0_st2_arr[12][7] <= 64'd18195737754871401302;
            ROM0_st2_arr[12][8] <= 64'd18446744060824649731;
            ROM0_st2_arr[12][9] <= 64'd2516679110167919243;
            ROM0_st2_arr[12][10] <= 64'd5354475383087621126;
            ROM0_st2_arr[12][11] <= 64'd7212304424746908984;
            ROM0_st2_arr[12][12] <= 64'd18446735273187346433;
            ROM0_st2_arr[12][13] <= 64'd4885406131420311944;
            ROM0_st2_arr[12][14] <= 64'd3183461194731576851;
            ROM0_st2_arr[12][15] <= 64'd15509998400778620264;
            ROM0_st2_arr[13][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[13][1] <= 64'd9818922367904463524;
            ROM0_st2_arr[13][2] <= 64'd151907467378121323;
            ROM0_st2_arr[13][3] <= 64'd14481943491905488994;
            ROM0_st2_arr[13][4] <= 64'd2251799813685256;
            ROM0_st2_arr[13][5] <= 64'd7159872751042635062;
            ROM0_st2_arr[13][6] <= 64'd14414733098329063675;
            ROM0_st2_arr[13][7] <= 64'd2189760912533326910;
            ROM0_st2_arr[13][8] <= 64'd576460752303423488;
            ROM0_st2_arr[13][9] <= 64'd8361668630589700543;
            ROM0_st2_arr[13][10] <= 64'd3739866984981691206;
            ROM0_st2_arr[13][11] <= 64'd5343314457212461663;
            ROM0_st2_arr[13][12] <= 64'd17179607036;
            ROM0_st2_arr[13][13] <= 64'd10192370097903824955;
            ROM0_st2_arr[13][14] <= 64'd3529731928842185170;
            ROM0_st2_arr[13][15] <= 64'd6578288040387767784;
            ROM0_st2_arr[14][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[14][1] <= 64'd822286005048470973;
            ROM0_st2_arr[14][2] <= 64'd9431669795342842913;
            ROM0_st2_arr[14][3] <= 64'd1633125474599800180;
            ROM0_st2_arr[14][4] <= 64'd281474976710655;
            ROM0_st2_arr[14][5] <= 64'd12787864249992692373;
            ROM0_st2_arr[14][6] <= 64'd17231484330389613737;
            ROM0_st2_arr[14][7] <= 64'd15858936941978258313;
            ROM0_st2_arr[14][8] <= 64'd18437736870159843329;
            ROM0_st2_arr[14][9] <= 64'd18328136608487584654;
            ROM0_st2_arr[14][10] <= 64'd6026834481055410692;
            ROM0_st2_arr[14][11] <= 64'd2966091928862697257;
            ROM0_st2_arr[14][12] <= 64'd144115188075856384;
            ROM0_st2_arr[14][13] <= 64'd5003087395582928323;
            ROM0_st2_arr[14][14] <= 64'd5079169390476357481;
            ROM0_st2_arr[14][15] <= 64'd12557198942430038686;
            ROM0_st2_arr[15][0] <= 64'd17293822565076172801;
            ROM0_st2_arr[15][1] <= 64'd7291801122603102867;
            ROM0_st2_arr[15][2] <= 64'd2391003455572333251;
            ROM0_st2_arr[15][3] <= 64'd5733718990552203475;
            ROM0_st2_arr[15][4] <= 64'd2305807824304734208;
            ROM0_st2_arr[15][5] <= 64'd17545206016321220698;
            ROM0_st2_arr[15][6] <= 64'd18314400042468094230;
            ROM0_st2_arr[15][7] <= 64'd15645300988549124365;
            ROM0_st2_arr[15][8] <= 64'd140737488355328;
            ROM0_st2_arr[15][9] <= 64'd611975439792384519;
            ROM0_st2_arr[15][10] <= 64'd18294836602036462998;
            ROM0_st2_arr[15][11] <= 64'd2229508537873380666;
            ROM0_st2_arr[15][12] <= 64'd18446462594437873666;
            ROM0_st2_arr[15][13] <= 64'd4764402665577370908;
            ROM0_st2_arr[15][14] <= 64'd1666382085084406020;
            ROM0_st2_arr[15][15] <= 64'd13493510495430156984;

            ROM0_st3_arr[0] <= 64'd17293822565076172801;
            ROM0_st3_arr[1] <= 64'd18014398505287680;
            ROM0_st3_arr[2] <= 64'd18446462594437939201;
            ROM0_st3_arr[3] <= 64'd4398046510080;
            ROM0_st3_arr[4] <= 64'd18446744000695107601;
            ROM0_st3_arr[5] <= 64'd4611686018427387904;
            ROM0_st3_arr[6] <= 64'd18374686475376656385;
            ROM0_st3_arr[7] <= 64'd1125899906842624;
            ROM0_st3_arr[8] <= 64'd18446726477228539905;
            ROM0_st3_arr[9] <= 64'd274877906944;
            ROM0_st3_arr[10] <= 64'd18446744065119617025;
            ROM0_st3_arr[11] <= 64'd67108864;
            ROM0_st3_arr[12] <= 64'd18446744069413535745;
            ROM0_st3_arr[13] <= 64'd16384;
            ROM0_st3_arr[14] <= 64'd18446744069414584065;
            ROM0_st3_arr[15] <= 64'd4;
            // ROM1 init
            ROM1_arr[0][0] <= 64'd1;
            ROM1_arr[0][1] <= 64'd1;
            ROM1_arr[0][2] <= 64'd1;
            ROM1_arr[0][3] <= 64'd1;
            ROM1_arr[0][4] <= 64'd1;
            ROM1_arr[0][5] <= 64'd1;
            ROM1_arr[0][6] <= 64'd1;
            ROM1_arr[0][7] <= 64'd1;
            ROM1_arr[0][8] <= 64'd1;
            ROM1_arr[0][9] <= 64'd1;
            ROM1_arr[0][10] <= 64'd1;
            ROM1_arr[0][11] <= 64'd1;
            ROM1_arr[0][12] <= 64'd1;
            ROM1_arr[0][13] <= 64'd1;
            ROM1_arr[0][14] <= 64'd1;
            ROM1_arr[0][15] <= 64'd1;
            ROM1_arr[1][0] <= 64'd1;
            ROM1_arr[1][1] <= 64'd17016677926152768545;
            ROM1_arr[1][2] <= 64'd2973809094719731252;
            ROM1_arr[1][3] <= 64'd8145372039058676274;
            ROM1_arr[1][4] <= 64'd6889485207579503204;
            ROM1_arr[1][5] <= 64'd453878597269088950;
            ROM1_arr[1][6] <= 64'd14799492472290523529;
            ROM1_arr[1][7] <= 64'd11526228256745639900;
            ROM1_arr[1][8] <= 64'd10006174791165856646;
            ROM1_arr[1][9] <= 64'd8463771714235575839;
            ROM1_arr[1][10] <= 64'd10450604126597135527;
            ROM1_arr[1][11] <= 64'd3953830850334785757;
            ROM1_arr[1][12] <= 64'd7190759909111520345;
            ROM1_arr[1][13] <= 64'd4619234339894857498;
            ROM1_arr[1][14] <= 64'd13250664030524184275;
            ROM1_arr[1][15] <= 64'd2180236998364722931;
            ROM1_arr[2][0] <= 64'd1;
            ROM1_arr[2][1] <= 64'd2973809094719731252;
            ROM1_arr[2][2] <= 64'd6889485207579503204;
            ROM1_arr[2][3] <= 64'd14799492472290523529;
            ROM1_arr[2][4] <= 64'd10006174791165856646;
            ROM1_arr[2][5] <= 64'd10450604126597135527;
            ROM1_arr[2][6] <= 64'd7190759909111520345;
            ROM1_arr[2][7] <= 64'd13250664030524184275;
            ROM1_arr[2][8] <= 64'd7059463857684370340;
            ROM1_arr[2][9] <= 64'd17011230650582925021;
            ROM1_arr[2][10] <= 64'd16905094363786184290;
            ROM1_arr[2][11] <= 64'd6238612790024380338;
            ROM1_arr[2][12] <= 64'd6702103175001071216;
            ROM1_arr[2][13] <= 64'd18208673802235871171;
            ROM1_arr[2][14] <= 64'd15984902507394762860;
            ROM1_arr[2][15] <= 64'd8445603439748857133;
            ROM1_arr[3][0] <= 64'd1;
            ROM1_arr[3][1] <= 64'd8145372039058676274;
            ROM1_arr[3][2] <= 64'd14799492472290523529;
            ROM1_arr[3][3] <= 64'd8463771714235575839;
            ROM1_arr[3][4] <= 64'd7190759909111520345;
            ROM1_arr[3][5] <= 64'd2180236998364722931;
            ROM1_arr[3][6] <= 64'd17011230650582925021;
            ROM1_arr[3][7] <= 64'd5770382478085514096;
            ROM1_arr[3][8] <= 64'd6702103175001071216;
            ROM1_arr[3][9] <= 64'd7650721134142770262;
            ROM1_arr[3][10] <= 64'd8445603439748857133;
            ROM1_arr[3][11] <= 64'd1633876473616625306;
            ROM1_arr[3][12] <= 64'd11102195893002206701;
            ROM1_arr[3][13] <= 64'd13030694632889454881;
            ROM1_arr[3][14] <= 64'd15253999561031414629;
            ROM1_arr[3][15] <= 64'd5194716592933687506;
            ROM1_arr[4][0] <= 64'd1;
            ROM1_arr[4][1] <= 64'd6889485207579503204;
            ROM1_arr[4][2] <= 64'd10006174791165856646;
            ROM1_arr[4][3] <= 64'd7190759909111520345;
            ROM1_arr[4][4] <= 64'd7059463857684370340;
            ROM1_arr[4][5] <= 64'd16905094363786184290;
            ROM1_arr[4][6] <= 64'd6702103175001071216;
            ROM1_arr[4][7] <= 64'd15984902507394762860;
            ROM1_arr[4][8] <= 64'd13835128420805115905;
            ROM1_arr[4][9] <= 64'd11102195893002206701;
            ROM1_arr[4][10] <= 64'd1897719374831994672;
            ROM1_arr[4][11] <= 64'd2128915576975457846;
            ROM1_arr[4][12] <= 64'd4442103655964903148;
            ROM1_arr[4][13] <= 64'd4156731661302306550;
            ROM1_arr[4][14] <= 64'd17920296056720464863;
            ROM1_arr[4][15] <= 64'd12365007338637617157;
            ROM1_arr[5][0] <= 64'd1;
            ROM1_arr[5][1] <= 64'd453878597269088950;
            ROM1_arr[5][2] <= 64'd10450604126597135527;
            ROM1_arr[5][3] <= 64'd2180236998364722931;
            ROM1_arr[5][4] <= 64'd16905094363786184290;
            ROM1_arr[5][5] <= 64'd642031755887803148;
            ROM1_arr[5][6] <= 64'd8445603439748857133;
            ROM1_arr[5][7] <= 64'd11384173023892451435;
            ROM1_arr[5][8] <= 64'd1897719374831994672;
            ROM1_arr[5][9] <= 64'd5194716592933687506;
            ROM1_arr[5][10] <= 64'd15908314874472904356;
            ROM1_arr[5][11] <= 64'd6212503712215198030;
            ROM1_arr[5][12] <= 64'd12365007338637617157;
            ROM1_arr[5][13] <= 64'd995696504716039625;
            ROM1_arr[5][14] <= 64'd9417275712919839734;
            ROM1_arr[5][15] <= 64'd14601330820526981151;
            ROM1_arr[6][0] <= 64'd1;
            ROM1_arr[6][1] <= 64'd14799492472290523529;
            ROM1_arr[6][2] <= 64'd7190759909111520345;
            ROM1_arr[6][3] <= 64'd17011230650582925021;
            ROM1_arr[6][4] <= 64'd6702103175001071216;
            ROM1_arr[6][5] <= 64'd8445603439748857133;
            ROM1_arr[6][6] <= 64'd11102195893002206701;
            ROM1_arr[6][7] <= 64'd15253999561031414629;
            ROM1_arr[6][8] <= 64'd4442103655964903148;
            ROM1_arr[6][9] <= 64'd13682879565831419937;
            ROM1_arr[6][10] <= 64'd12365007338637617157;
            ROM1_arr[6][11] <= 64'd12806605743856568005;
            ROM1_arr[6][12] <= 64'd13533145890581203496;
            ROM1_arr[6][13] <= 64'd10156112135473104598;
            ROM1_arr[6][14] <= 64'd4576915052531526319;
            ROM1_arr[6][15] <= 64'd11998590678972281283;
            ROM1_arr[7][0] <= 64'd1;
            ROM1_arr[7][1] <= 64'd11526228256745639900;
            ROM1_arr[7][2] <= 64'd13250664030524184275;
            ROM1_arr[7][3] <= 64'd5770382478085514096;
            ROM1_arr[7][4] <= 64'd15984902507394762860;
            ROM1_arr[7][5] <= 64'd11384173023892451435;
            ROM1_arr[7][6] <= 64'd15253999561031414629;
            ROM1_arr[7][7] <= 64'd16251565245213924195;
            ROM1_arr[7][8] <= 64'd17920296056720464863;
            ROM1_arr[7][9] <= 64'd5004020984668548385;
            ROM1_arr[7][10] <= 64'd9417275712919839734;
            ROM1_arr[7][11] <= 64'd6631640021333632646;
            ROM1_arr[7][12] <= 64'd4576915052531526319;
            ROM1_arr[7][13] <= 64'd9499642494161596470;
            ROM1_arr[7][14] <= 64'd10026248927784619520;
            ROM1_arr[7][15] <= 64'd13015839270796764972;
            ROM1_arr[8][0] <= 64'd1;
            ROM1_arr[8][1] <= 64'd10006174791165856646;
            ROM1_arr[8][2] <= 64'd7059463857684370340;
            ROM1_arr[8][3] <= 64'd6702103175001071216;
            ROM1_arr[8][4] <= 64'd13835128420805115905;
            ROM1_arr[8][5] <= 64'd1897719374831994672;
            ROM1_arr[8][6] <= 64'd4442103655964903148;
            ROM1_arr[8][7] <= 64'd17920296056720464863;
            ROM1_arr[8][8] <= 64'd35184372088832;
            ROM1_arr[8][9] <= 64'd13533145890581203496;
            ROM1_arr[8][10] <= 64'd10561990880479197442;
            ROM1_arr[8][11] <= 64'd17345757166192390690;
            ROM1_arr[8][12] <= 64'd576469548262227968;
            ROM1_arr[8][13] <= 64'd6529358023436602414;
            ROM1_arr[8][14] <= 64'd13949104517951277988;
            ROM1_arr[8][15] <= 64'd4126998567329314197;
            ROM1_arr[9][0] <= 64'd1;
            ROM1_arr[9][1] <= 64'd8463771714235575839;
            ROM1_arr[9][2] <= 64'd17011230650582925021;
            ROM1_arr[9][3] <= 64'd7650721134142770262;
            ROM1_arr[9][4] <= 64'd11102195893002206701;
            ROM1_arr[9][5] <= 64'd5194716592933687506;
            ROM1_arr[9][6] <= 64'd13682879565831419937;
            ROM1_arr[9][7] <= 64'd5004020984668548385;
            ROM1_arr[9][8] <= 64'd13533145890581203496;
            ROM1_arr[9][9] <= 64'd11050185740979045171;
            ROM1_arr[9][10] <= 64'd11998590678972281283;
            ROM1_arr[9][11] <= 64'd14748993927606327403;
            ROM1_arr[9][12] <= 64'd14804671509201811970;
            ROM1_arr[9][13] <= 64'd9853084201154921057;
            ROM1_arr[9][14] <= 64'd7835252777128489741;
            ROM1_arr[9][15] <= 64'd7890353213857230017;
            ROM1_arr[10][0] <= 64'd1;
            ROM1_arr[10][1] <= 64'd10450604126597135527;
            ROM1_arr[10][2] <= 64'd16905094363786184290;
            ROM1_arr[10][3] <= 64'd8445603439748857133;
            ROM1_arr[10][4] <= 64'd1897719374831994672;
            ROM1_arr[10][5] <= 64'd15908314874472904356;
            ROM1_arr[10][6] <= 64'd12365007338637617157;
            ROM1_arr[10][7] <= 64'd9417275712919839734;
            ROM1_arr[10][8] <= 64'd10561990880479197442;
            ROM1_arr[10][9] <= 64'd11998590678972281283;
            ROM1_arr[10][10] <= 64'd12486396704535672088;
            ROM1_arr[10][11] <= 64'd3854327039422012671;
            ROM1_arr[10][12] <= 64'd4126998567329314197;
            ROM1_arr[10][13] <= 64'd14941513789294353960;
            ROM1_arr[10][14] <= 64'd7093403778535204495;
            ROM1_arr[10][15] <= 64'd14314040479386013058;
            ROM1_arr[11][0] <= 64'd1;
            ROM1_arr[11][1] <= 64'd3953830850334785757;
            ROM1_arr[11][2] <= 64'd6238612790024380338;
            ROM1_arr[11][3] <= 64'd1633876473616625306;
            ROM1_arr[11][4] <= 64'd2128915576975457846;
            ROM1_arr[11][5] <= 64'd6212503712215198030;
            ROM1_arr[11][6] <= 64'd12806605743856568005;
            ROM1_arr[11][7] <= 64'd6631640021333632646;
            ROM1_arr[11][8] <= 64'd17345757166192390690;
            ROM1_arr[11][9] <= 64'd14748993927606327403;
            ROM1_arr[11][10] <= 64'd3854327039422012671;
            ROM1_arr[11][11] <= 64'd6572141765742720031;
            ROM1_arr[11][12] <= 64'd10268645332677273943;
            ROM1_arr[11][13] <= 64'd14665682977215298085;
            ROM1_arr[11][14] <= 64'd580180600093873153;
            ROM1_arr[11][15] <= 64'd652687206561795469;
            ROM1_arr[12][0] <= 64'd1;
            ROM1_arr[12][1] <= 64'd7190759909111520345;
            ROM1_arr[12][2] <= 64'd6702103175001071216;
            ROM1_arr[12][3] <= 64'd11102195893002206701;
            ROM1_arr[12][4] <= 64'd4442103655964903148;
            ROM1_arr[12][5] <= 64'd12365007338637617157;
            ROM1_arr[12][6] <= 64'd13533145890581203496;
            ROM1_arr[12][7] <= 64'd4576915052531526319;
            ROM1_arr[12][8] <= 64'd576469548262227968;
            ROM1_arr[12][9] <= 64'd14804671509201811970;
            ROM1_arr[12][10] <= 64'd4126998567329314197;
            ROM1_arr[12][11] <= 64'd10268645332677273943;
            ROM1_arr[12][12] <= 64'd10265989416269385394;
            ROM1_arr[12][13] <= 64'd12432372446044483551;
            ROM1_arr[12][14] <= 64'd13805406186829188324;
            ROM1_arr[12][15] <= 64'd15499491376360706981;
            ROM1_arr[13][0] <= 64'd1;
            ROM1_arr[13][1] <= 64'd4619234339894857498;
            ROM1_arr[13][2] <= 64'd18208673802235871171;
            ROM1_arr[13][3] <= 64'd13030694632889454881;
            ROM1_arr[13][4] <= 64'd4156731661302306550;
            ROM1_arr[13][5] <= 64'd995696504716039625;
            ROM1_arr[13][6] <= 64'd10156112135473104598;
            ROM1_arr[13][7] <= 64'd9499642494161596470;
            ROM1_arr[13][8] <= 64'd6529358023436602414;
            ROM1_arr[13][9] <= 64'd9853084201154921057;
            ROM1_arr[13][10] <= 64'd14941513789294353960;
            ROM1_arr[13][11] <= 64'd14665682977215298085;
            ROM1_arr[13][12] <= 64'd12432372446044483551;
            ROM1_arr[13][13] <= 64'd11997839738651575743;
            ROM1_arr[13][14] <= 64'd9297807417575779104;
            ROM1_arr[13][15] <= 64'd13545855348012112781;
            ROM1_arr[14][0] <= 64'd1;
            ROM1_arr[14][1] <= 64'd13250664030524184275;
            ROM1_arr[14][2] <= 64'd15984902507394762860;
            ROM1_arr[14][3] <= 64'd15253999561031414629;
            ROM1_arr[14][4] <= 64'd17920296056720464863;
            ROM1_arr[14][5] <= 64'd9417275712919839734;
            ROM1_arr[14][6] <= 64'd4576915052531526319;
            ROM1_arr[14][7] <= 64'd10026248927784619520;
            ROM1_arr[14][8] <= 64'd13949104517951277988;
            ROM1_arr[14][9] <= 64'd7835252777128489741;
            ROM1_arr[14][10] <= 64'd7093403778535204495;
            ROM1_arr[14][11] <= 64'd580180600093873153;
            ROM1_arr[14][12] <= 64'd13805406186829188324;
            ROM1_arr[14][13] <= 64'd9297807417575779104;
            ROM1_arr[14][14] <= 64'd12032395915935294938;
            ROM1_arr[14][15] <= 64'd15581468049507881811;
            ROM1_arr[15][0] <= 64'd1;
            ROM1_arr[15][1] <= 64'd2180236998364722931;
            ROM1_arr[15][2] <= 64'd8445603439748857133;
            ROM1_arr[15][3] <= 64'd5194716592933687506;
            ROM1_arr[15][4] <= 64'd12365007338637617157;
            ROM1_arr[15][5] <= 64'd14601330820526981151;
            ROM1_arr[15][6] <= 64'd11998590678972281283;
            ROM1_arr[15][7] <= 64'd13015839270796764972;
            ROM1_arr[15][8] <= 64'd4126998567329314197;
            ROM1_arr[15][9] <= 64'd7890353213857230017;
            ROM1_arr[15][10] <= 64'd14314040479386013058;
            ROM1_arr[15][11] <= 64'd652687206561795469;
            ROM1_arr[15][12] <= 64'd15499491376360706981;
            ROM1_arr[15][13] <= 64'd13545855348012112781;
            ROM1_arr[15][14] <= 64'd15581468049507881811;
            ROM1_arr[15][15] <= 64'd4967386273503838092;
            // ROM2 init
            ROM2_arr[0][0] <= 64'd1;
            ROM2_arr[0][1] <= 64'd1;
            ROM2_arr[0][2] <= 64'd1;
            ROM2_arr[0][3] <= 64'd1;
            ROM2_arr[0][4] <= 64'd1;
            ROM2_arr[0][5] <= 64'd1;
            ROM2_arr[0][6] <= 64'd1;
            ROM2_arr[0][7] <= 64'd1;
            ROM2_arr[0][8] <= 64'd1;
            ROM2_arr[0][9] <= 64'd1;
            ROM2_arr[0][10] <= 64'd1;
            ROM2_arr[0][11] <= 64'd1;
            ROM2_arr[0][12] <= 64'd1;
            ROM2_arr[0][13] <= 64'd1;
            ROM2_arr[0][14] <= 64'd1;
            ROM2_arr[0][15] <= 64'd1;
            ROM2_arr[1][0] <= 64'd1;
            ROM2_arr[1][1] <= 64'd8442954237739851301;
            ROM2_arr[1][2] <= 64'd8296420140406050866;
            ROM2_arr[1][3] <= 64'd8975318665775642004;
            ROM2_arr[1][4] <= 64'd14570053890742115847;
            ROM2_arr[1][5] <= 64'd9712494135743485235;
            ROM2_arr[1][6] <= 64'd8520458930592089940;
            ROM2_arr[1][7] <= 64'd5442418197918194943;
            ROM2_arr[1][8] <= 64'd459643346215618215;
            ROM2_arr[1][9] <= 64'd8477580977336904871;
            ROM2_arr[1][10] <= 64'd2571862908476870164;
            ROM2_arr[1][11] <= 64'd730718612094303599;
            ROM2_arr[1][12] <= 64'd16027583595078457158;
            ROM2_arr[1][13] <= 64'd15790091985445428011;
            ROM2_arr[1][14] <= 64'd15636908079422696657;
            ROM2_arr[1][15] <= 64'd14500624711942570790;
            ROM2_arr[2][0] <= 64'd1;
            ROM2_arr[2][1] <= 64'd8296420140406050866;
            ROM2_arr[2][2] <= 64'd14570053890742115847;
            ROM2_arr[2][3] <= 64'd8520458930592089940;
            ROM2_arr[2][4] <= 64'd459643346215618215;
            ROM2_arr[2][5] <= 64'd2571862908476870164;
            ROM2_arr[2][6] <= 64'd16027583595078457158;
            ROM2_arr[2][7] <= 64'd15636908079422696657;
            ROM2_arr[2][8] <= 64'd17016677926152768545;
            ROM2_arr[2][9] <= 64'd15354180691825273826;
            ROM2_arr[2][10] <= 64'd2642934261869995837;
            ROM2_arr[2][11] <= 64'd12120845767179702978;
            ROM2_arr[2][12] <= 64'd9704267196562286842;
            ROM2_arr[2][13] <= 64'd8303301787244588674;
            ROM2_arr[2][14] <= 64'd15097984348022460756;
            ROM2_arr[2][15] <= 64'd9254204077078059724;
            ROM2_arr[3][0] <= 64'd1;
            ROM2_arr[3][1] <= 64'd8975318665775642004;
            ROM2_arr[3][2] <= 64'd8520458930592089940;
            ROM2_arr[3][3] <= 64'd8477580977336904871;
            ROM2_arr[3][4] <= 64'd16027583595078457158;
            ROM2_arr[3][5] <= 64'd14500624711942570790;
            ROM2_arr[3][6] <= 64'd15354180691825273826;
            ROM2_arr[3][7] <= 64'd14123590475017358834;
            ROM2_arr[3][8] <= 64'd9704267196562286842;
            ROM2_arr[3][9] <= 64'd17759015114171266566;
            ROM2_arr[3][10] <= 64'd9254204077078059724;
            ROM2_arr[3][11] <= 64'd3502348020251649926;
            ROM2_arr[3][12] <= 64'd3634574816773780305;
            ROM2_arr[3][13] <= 64'd5597741650023885745;
            ROM2_arr[3][14] <= 64'd12860603398506203576;
            ROM2_arr[3][15] <= 64'd6088724424422443500;
            ROM2_arr[4][0] <= 64'd1;
            ROM2_arr[4][1] <= 64'd14570053890742115847;
            ROM2_arr[4][2] <= 64'd459643346215618215;
            ROM2_arr[4][3] <= 64'd16027583595078457158;
            ROM2_arr[4][4] <= 64'd17016677926152768545;
            ROM2_arr[4][5] <= 64'd2642934261869995837;
            ROM2_arr[4][6] <= 64'd9704267196562286842;
            ROM2_arr[4][7] <= 64'd15097984348022460756;
            ROM2_arr[4][8] <= 64'd2973809094719731252;
            ROM2_arr[4][9] <= 64'd3634574816773780305;
            ROM2_arr[4][10] <= 64'd17738676007726690413;
            ROM2_arr[4][11] <= 64'd9105921508417528907;
            ROM2_arr[4][12] <= 64'd8145372039058676274;
            ROM2_arr[4][13] <= 64'd13284953271058402611;
            ROM2_arr[4][14] <= 64'd7937777424398523163;
            ROM2_arr[4][15] <= 64'd8925204892929839437;
            ROM2_arr[5][0] <= 64'd1;
            ROM2_arr[5][1] <= 64'd9712494135743485235;
            ROM2_arr[5][2] <= 64'd2571862908476870164;
            ROM2_arr[5][3] <= 64'd14500624711942570790;
            ROM2_arr[5][4] <= 64'd2642934261869995837;
            ROM2_arr[5][5] <= 64'd13177409762334527172;
            ROM2_arr[5][6] <= 64'd9254204077078059724;
            ROM2_arr[5][7] <= 64'd18310129038502196404;
            ROM2_arr[5][8] <= 64'd17738676007726690413;
            ROM2_arr[5][9] <= 64'd6088724424422443500;
            ROM2_arr[5][10] <= 64'd2064229586559886558;
            ROM2_arr[5][11] <= 64'd10529815446215197801;
            ROM2_arr[5][12] <= 64'd8925204892929839437;
            ROM2_arr[5][13] <= 64'd7251235515904981255;
            ROM2_arr[5][14] <= 64'd6072555943748209899;
            ROM2_arr[5][15] <= 64'd1741246929451345145;
            ROM2_arr[6][0] <= 64'd1;
            ROM2_arr[6][1] <= 64'd8520458930592089940;
            ROM2_arr[6][2] <= 64'd16027583595078457158;
            ROM2_arr[6][3] <= 64'd15354180691825273826;
            ROM2_arr[6][4] <= 64'd9704267196562286842;
            ROM2_arr[6][5] <= 64'd9254204077078059724;
            ROM2_arr[6][6] <= 64'd3634574816773780305;
            ROM2_arr[6][7] <= 64'd12860603398506203576;
            ROM2_arr[6][8] <= 64'd8145372039058676274;
            ROM2_arr[6][9] <= 64'd17924415806212830485;
            ROM2_arr[6][10] <= 64'd8925204892929839437;
            ROM2_arr[6][11] <= 64'd1369635493243148371;
            ROM2_arr[6][12] <= 64'd16843210144819986575;
            ROM2_arr[6][13] <= 64'd9324490876611876183;
            ROM2_arr[6][14] <= 64'd11511052703523625381;
            ROM2_arr[6][15] <= 64'd3657254226843515683;
            ROM2_arr[7][0] <= 64'd1;
            ROM2_arr[7][1] <= 64'd5442418197918194943;
            ROM2_arr[7][2] <= 64'd15636908079422696657;
            ROM2_arr[7][3] <= 64'd14123590475017358834;
            ROM2_arr[7][4] <= 64'd15097984348022460756;
            ROM2_arr[7][5] <= 64'd18310129038502196404;
            ROM2_arr[7][6] <= 64'd12860603398506203576;
            ROM2_arr[7][7] <= 64'd2928469370849851995;
            ROM2_arr[7][8] <= 64'd7937777424398523163;
            ROM2_arr[7][9] <= 64'd9111473011521032935;
            ROM2_arr[7][10] <= 64'd6072555943748209899;
            ROM2_arr[7][11] <= 64'd17589514971603809675;
            ROM2_arr[7][12] <= 64'd11511052703523625381;
            ROM2_arr[7][13] <= 64'd4131273418538853697;
            ROM2_arr[7][14] <= 64'd9725369440298319348;
            ROM2_arr[7][15] <= 64'd8026948575168308684;
            ROM2_arr[8][0] <= 64'd1;
            ROM2_arr[8][1] <= 64'd459643346215618215;
            ROM2_arr[8][2] <= 64'd17016677926152768545;
            ROM2_arr[8][3] <= 64'd9704267196562286842;
            ROM2_arr[8][4] <= 64'd2973809094719731252;
            ROM2_arr[8][5] <= 64'd17738676007726690413;
            ROM2_arr[8][6] <= 64'd8145372039058676274;
            ROM2_arr[8][7] <= 64'd7937777424398523163;
            ROM2_arr[8][8] <= 64'd6889485207579503204;
            ROM2_arr[8][9] <= 64'd16843210144819986575;
            ROM2_arr[8][10] <= 64'd453878597269088950;
            ROM2_arr[8][11] <= 64'd1944587153055514591;
            ROM2_arr[8][12] <= 64'd14799492472290523529;
            ROM2_arr[8][13] <= 64'd5546020403660220517;
            ROM2_arr[8][14] <= 64'd11526228256745639900;
            ROM2_arr[8][15] <= 64'd7583194663533335603;
            ROM2_arr[9][0] <= 64'd1;
            ROM2_arr[9][1] <= 64'd8477580977336904871;
            ROM2_arr[9][2] <= 64'd15354180691825273826;
            ROM2_arr[9][3] <= 64'd17759015114171266566;
            ROM2_arr[9][4] <= 64'd3634574816773780305;
            ROM2_arr[9][5] <= 64'd6088724424422443500;
            ROM2_arr[9][6] <= 64'd17924415806212830485;
            ROM2_arr[9][7] <= 64'd9111473011521032935;
            ROM2_arr[9][8] <= 64'd16843210144819986575;
            ROM2_arr[9][9] <= 64'd3001722651578882312;
            ROM2_arr[9][10] <= 64'd3657254226843515683;
            ROM2_arr[9][11] <= 64'd5325893774437366420;
            ROM2_arr[9][12] <= 64'd12671531405601353448;
            ROM2_arr[9][13] <= 64'd3032592923511514202;
            ROM2_arr[9][14] <= 64'd9792896423618660571;
            ROM2_arr[9][15] <= 64'd12622989934929842507;
            ROM2_arr[10][0] <= 64'd1;
            ROM2_arr[10][1] <= 64'd2571862908476870164;
            ROM2_arr[10][2] <= 64'd2642934261869995837;
            ROM2_arr[10][3] <= 64'd9254204077078059724;
            ROM2_arr[10][4] <= 64'd17738676007726690413;
            ROM2_arr[10][5] <= 64'd2064229586559886558;
            ROM2_arr[10][6] <= 64'd8925204892929839437;
            ROM2_arr[10][7] <= 64'd6072555943748209899;
            ROM2_arr[10][8] <= 64'd453878597269088950;
            ROM2_arr[10][9] <= 64'd3657254226843515683;
            ROM2_arr[10][10] <= 64'd9044778990070702823;
            ROM2_arr[10][11] <= 64'd12748278382855927485;
            ROM2_arr[10][12] <= 64'd7583194663533335603;
            ROM2_arr[10][13] <= 64'd17697369196786003250;
            ROM2_arr[10][14] <= 64'd15686100554272703417;
            ROM2_arr[10][15] <= 64'd17323211596453562164;
            ROM2_arr[11][0] <= 64'd1;
            ROM2_arr[11][1] <= 64'd730718612094303599;
            ROM2_arr[11][2] <= 64'd12120845767179702978;
            ROM2_arr[11][3] <= 64'd3502348020251649926;
            ROM2_arr[11][4] <= 64'd9105921508417528907;
            ROM2_arr[11][5] <= 64'd10529815446215197801;
            ROM2_arr[11][6] <= 64'd1369635493243148371;
            ROM2_arr[11][7] <= 64'd17589514971603809675;
            ROM2_arr[11][8] <= 64'd1944587153055514591;
            ROM2_arr[11][9] <= 64'd5325893774437366420;
            ROM2_arr[11][10] <= 64'd12748278382855927485;
            ROM2_arr[11][11] <= 64'd14075137670294329533;
            ROM2_arr[11][12] <= 64'd17165287979911939135;
            ROM2_arr[11][13] <= 64'd16015250250966057106;
            ROM2_arr[11][14] <= 64'd17793898918920342346;
            ROM2_arr[11][15] <= 64'd14059751200357075018;
            ROM2_arr[12][0] <= 64'd1;
            ROM2_arr[12][1] <= 64'd16027583595078457158;
            ROM2_arr[12][2] <= 64'd9704267196562286842;
            ROM2_arr[12][3] <= 64'd3634574816773780305;
            ROM2_arr[12][4] <= 64'd8145372039058676274;
            ROM2_arr[12][5] <= 64'd8925204892929839437;
            ROM2_arr[12][6] <= 64'd16843210144819986575;
            ROM2_arr[12][7] <= 64'd11511052703523625381;
            ROM2_arr[12][8] <= 64'd14799492472290523529;
            ROM2_arr[12][9] <= 64'd12671531405601353448;
            ROM2_arr[12][10] <= 64'd7583194663533335603;
            ROM2_arr[12][11] <= 64'd17165287979911939135;
            ROM2_arr[12][12] <= 64'd8463771714235575839;
            ROM2_arr[12][13] <= 64'd13304357142560244146;
            ROM2_arr[12][14] <= 64'd6743138205473560756;
            ROM2_arr[12][15] <= 64'd16372052743821334332;
            ROM2_arr[13][0] <= 64'd1;
            ROM2_arr[13][1] <= 64'd15790091985445428011;
            ROM2_arr[13][2] <= 64'd8303301787244588674;
            ROM2_arr[13][3] <= 64'd5597741650023885745;
            ROM2_arr[13][4] <= 64'd13284953271058402611;
            ROM2_arr[13][5] <= 64'd7251235515904981255;
            ROM2_arr[13][6] <= 64'd9324490876611876183;
            ROM2_arr[13][7] <= 64'd4131273418538853697;
            ROM2_arr[13][8] <= 64'd5546020403660220517;
            ROM2_arr[13][9] <= 64'd3032592923511514202;
            ROM2_arr[13][10] <= 64'd17697369196786003250;
            ROM2_arr[13][11] <= 64'd16015250250966057106;
            ROM2_arr[13][12] <= 64'd13304357142560244146;
            ROM2_arr[13][13] <= 64'd855610743119371585;
            ROM2_arr[13][14] <= 64'd18262221851015199223;
            ROM2_arr[13][15] <= 64'd10989941768648740935;
            ROM2_arr[14][0] <= 64'd1;
            ROM2_arr[14][1] <= 64'd15636908079422696657;
            ROM2_arr[14][2] <= 64'd15097984348022460756;
            ROM2_arr[14][3] <= 64'd12860603398506203576;
            ROM2_arr[14][4] <= 64'd7937777424398523163;
            ROM2_arr[14][5] <= 64'd6072555943748209899;
            ROM2_arr[14][6] <= 64'd11511052703523625381;
            ROM2_arr[14][7] <= 64'd9725369440298319348;
            ROM2_arr[14][8] <= 64'd11526228256745639900;
            ROM2_arr[14][9] <= 64'd9792896423618660571;
            ROM2_arr[14][10] <= 64'd15686100554272703417;
            ROM2_arr[14][11] <= 64'd17793898918920342346;
            ROM2_arr[14][12] <= 64'd6743138205473560756;
            ROM2_arr[14][13] <= 64'd18262221851015199223;
            ROM2_arr[14][14] <= 64'd10542535943374472194;
            ROM2_arr[14][15] <= 64'd8468994490826810714;
            ROM2_arr[15][0] <= 64'd1;
            ROM2_arr[15][1] <= 64'd14500624711942570790;
            ROM2_arr[15][2] <= 64'd9254204077078059724;
            ROM2_arr[15][3] <= 64'd6088724424422443500;
            ROM2_arr[15][4] <= 64'd8925204892929839437;
            ROM2_arr[15][5] <= 64'd1741246929451345145;
            ROM2_arr[15][6] <= 64'd3657254226843515683;
            ROM2_arr[15][7] <= 64'd8026948575168308684;
            ROM2_arr[15][8] <= 64'd7583194663533335603;
            ROM2_arr[15][9] <= 64'd12622989934929842507;
            ROM2_arr[15][10] <= 64'd17323211596453562164;
            ROM2_arr[15][11] <= 64'd14059751200357075018;
            ROM2_arr[15][12] <= 64'd16372052743821334332;
            ROM2_arr[15][13] <= 64'd10989941768648740935;
            ROM2_arr[15][14] <= 64'd8468994490826810714;
            ROM2_arr[15][15] <= 64'd5457663874430016353;
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM0_b0     <= 64'd0    ;
            ROM0_b1     <= 64'd0    ;
            ROM0_b2     <= 64'd0    ;
            ROM0_b3     <= 64'd0    ;
            ROM0_b4     <= 64'd0    ;
            ROM0_b5     <= 64'd0    ;
            ROM0_b6     <= 64'd0    ;
            ROM0_b7     <= 64'd0    ;
            ROM0_b8     <= 64'd0    ;
            ROM0_b9     <= 64'd0    ;
            ROM0_b10    <= 64'd0    ;
            ROM0_b11    <= 64'd0    ;
            ROM0_b12    <= 64'd0    ; 
            ROM0_b13    <= 64'd0    ;
            ROM0_b14    <= 64'd0    ; 
            ROM0_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (FFT_stage_in)
                    2'd0: begin
                        case (MA0)
                            4'd0:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[0][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[0][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[0][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[0][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[0][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[0][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[0][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[0][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[0][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[0][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[0][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[0][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[0][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[0][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[0][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[0][15] ;
                                end
                            4'd1:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[1][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[1][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[1][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[1][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[1][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[1][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[1][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[1][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[1][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[1][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[1][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[1][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[1][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[1][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[1][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[1][15] ;
                                end
                            4'd2:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[2][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[2][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[2][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[2][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[2][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[2][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[2][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[2][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[2][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[2][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[2][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[2][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[2][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[2][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[2][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[2][15] ;
                                end
                            4'd3:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[3][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[3][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[3][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[3][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[3][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[3][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[3][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[3][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[3][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[3][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[3][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[3][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[3][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[3][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[3][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[3][15] ;
                                end
                            4'd4:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[4][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[4][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[4][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[4][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[4][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[4][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[4][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[4][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[4][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[4][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[4][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[4][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[4][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[4][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[4][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[4][15] ;
                                end
                            4'd5:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[5][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[5][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[5][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[5][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[5][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[5][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[5][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[5][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[5][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[5][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[5][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[5][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[5][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[5][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[5][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[5][15] ;
                                end
                            4'd6:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[6][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[6][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[6][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[6][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[6][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[6][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[6][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[6][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[6][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[6][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[6][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[6][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[6][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[6][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[6][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[6][15] ;
                                end
                            4'd7:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[7][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[7][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[7][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[7][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[7][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[7][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[7][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[7][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[7][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[7][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[7][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[7][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[7][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[7][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[7][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[7][15] ;
                                end
                            4'd8:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[8][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[8][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[8][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[8][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[8][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[8][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[8][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[8][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[8][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[8][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[8][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[8][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[8][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[8][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[8][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[8][15] ;
                                end
                            4'd9:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[9][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[9][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[9][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[9][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[9][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[9][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[9][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[9][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[9][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[9][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[9][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[9][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[9][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[9][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[9][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[9][15] ;
                                end
                            4'd10:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[10][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[10][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[10][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[10][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[10][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[10][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[10][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[10][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[10][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[10][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[10][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[10][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[10][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[10][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[10][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[10][15] ;
                                end
                            4'd11:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[11][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[11][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[11][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[11][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[11][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[11][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[11][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[11][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[11][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[11][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[11][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[11][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[11][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[11][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[11][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[11][15] ;
                                end
                            4'd12:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[12][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[12][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[12][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[12][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[12][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[12][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[12][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[12][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[12][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[12][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[12][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[12][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[12][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[12][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[12][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[12][15] ;
                                end
                            4'd13:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[13][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[13][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[13][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[13][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[13][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[13][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[13][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[13][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[13][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[13][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[13][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[13][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[13][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[13][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[13][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[13][15] ;
                                end
                            4'd14:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[14][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[14][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[14][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[14][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[14][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[14][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[14][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[14][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[14][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[14][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[14][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[14][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[14][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[14][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[14][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[14][15] ;
                                end
                            4'd15:
                                begin
                                    ROM0_b0     <=  ROM0_st0_arr[15][0]  ;
                                    ROM0_b1     <=  ROM0_st0_arr[15][1]  ;
                                    ROM0_b2     <=  ROM0_st0_arr[15][2]  ;
                                    ROM0_b3     <=  ROM0_st0_arr[15][3]  ;
                                    ROM0_b4     <=  ROM0_st0_arr[15][4]  ;
                                    ROM0_b5     <=  ROM0_st0_arr[15][5]  ;
                                    ROM0_b6     <=  ROM0_st0_arr[15][6]  ;
                                    ROM0_b7     <=  ROM0_st0_arr[15][7]  ;
                                    ROM0_b8     <=  ROM0_st0_arr[15][8]  ;
                                    ROM0_b9     <=  ROM0_st0_arr[15][9]  ;
                                    ROM0_b10    <=  ROM0_st0_arr[15][10] ;
                                    ROM0_b11    <=  ROM0_st0_arr[15][11] ;
                                    ROM0_b12    <=  ROM0_st0_arr[15][12] ;
                                    ROM0_b13    <=  ROM0_st0_arr[15][13] ;
                                    ROM0_b14    <=  ROM0_st0_arr[15][14] ;
                                    ROM0_b15    <=  ROM0_st0_arr[15][15] ;
                                end
                        endcase
                    end
                    2'd1: begin
                        case (MA0)
                            4'd0:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[0][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[0][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[0][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[0][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[0][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[0][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[0][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[0][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[0][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[0][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[0][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[0][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[0][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[0][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[0][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[0][15] ;
                                end
                            4'd1:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[1][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[1][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[1][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[1][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[1][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[1][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[1][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[1][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[1][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[1][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[1][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[1][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[1][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[1][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[1][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[1][15] ;
                                end
                            4'd2:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[2][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[2][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[2][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[2][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[2][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[2][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[2][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[2][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[2][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[2][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[2][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[2][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[2][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[2][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[2][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[2][15] ;
                                end
                            4'd3:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[3][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[3][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[3][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[3][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[3][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[3][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[3][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[3][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[3][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[3][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[3][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[3][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[3][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[3][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[3][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[3][15] ;
                                end
                            4'd4:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[4][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[4][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[4][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[4][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[4][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[4][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[4][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[4][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[4][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[4][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[4][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[4][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[4][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[4][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[4][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[4][15] ;
                                end
                            4'd5:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[5][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[5][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[5][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[5][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[5][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[5][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[5][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[5][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[5][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[5][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[5][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[5][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[5][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[5][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[5][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[5][15] ;
                                end
                            4'd6:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[6][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[6][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[6][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[6][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[6][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[6][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[6][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[6][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[6][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[6][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[6][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[6][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[6][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[6][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[6][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[6][15] ;
                                end
                            4'd7:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[7][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[7][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[7][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[7][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[7][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[7][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[7][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[7][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[7][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[7][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[7][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[7][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[7][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[7][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[7][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[7][15] ;
                                end
                            4'd8:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[8][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[8][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[8][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[8][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[8][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[8][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[8][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[8][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[8][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[8][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[8][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[8][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[8][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[8][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[8][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[8][15] ;
                                end
                            4'd9:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[9][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[9][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[9][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[9][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[9][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[9][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[9][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[9][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[9][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[9][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[9][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[9][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[9][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[9][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[9][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[9][15] ;
                                end
                            4'd10:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[10][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[10][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[10][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[10][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[10][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[10][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[10][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[10][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[10][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[10][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[10][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[10][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[10][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[10][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[10][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[10][15] ;
                                end
                            4'd11:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[11][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[11][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[11][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[11][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[11][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[11][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[11][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[11][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[11][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[11][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[11][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[11][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[11][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[11][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[11][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[11][15] ;
                                end
                            4'd12:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[12][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[12][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[12][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[12][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[12][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[12][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[12][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[12][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[12][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[12][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[12][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[12][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[12][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[12][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[12][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[12][15] ;
                                end
                            4'd13:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[13][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[13][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[13][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[13][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[13][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[13][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[13][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[13][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[13][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[13][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[13][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[13][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[13][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[13][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[13][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[13][15] ;
                                end
                            4'd14:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[14][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[14][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[14][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[14][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[14][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[14][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[14][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[14][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[14][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[14][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[14][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[14][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[14][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[14][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[14][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[14][15] ;
                                end
                            4'd15:
                                begin
                                    ROM0_b0     <=  ROM0_st1_arr[15][0]  ;
                                    ROM0_b1     <=  ROM0_st1_arr[15][1]  ;
                                    ROM0_b2     <=  ROM0_st1_arr[15][2]  ;
                                    ROM0_b3     <=  ROM0_st1_arr[15][3]  ;
                                    ROM0_b4     <=  ROM0_st1_arr[15][4]  ;
                                    ROM0_b5     <=  ROM0_st1_arr[15][5]  ;
                                    ROM0_b6     <=  ROM0_st1_arr[15][6]  ;
                                    ROM0_b7     <=  ROM0_st1_arr[15][7]  ;
                                    ROM0_b8     <=  ROM0_st1_arr[15][8]  ;
                                    ROM0_b9     <=  ROM0_st1_arr[15][9]  ;
                                    ROM0_b10    <=  ROM0_st1_arr[15][10] ;
                                    ROM0_b11    <=  ROM0_st1_arr[15][11] ;
                                    ROM0_b12    <=  ROM0_st1_arr[15][12] ;
                                    ROM0_b13    <=  ROM0_st1_arr[15][13] ;
                                    ROM0_b14    <=  ROM0_st1_arr[15][14] ;
                                    ROM0_b15    <=  ROM0_st1_arr[15][15] ;
                                end
                        endcase
                    end
                    2'd2: begin
                        case (MA0)
                            4'd0:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[0][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[0][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[0][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[0][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[0][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[0][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[0][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[0][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[0][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[0][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[0][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[0][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[0][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[0][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[0][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[0][15] ;
                                end
                            4'd1:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[1][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[1][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[1][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[1][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[1][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[1][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[1][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[1][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[1][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[1][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[1][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[1][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[1][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[1][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[1][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[1][15] ;
                                end
                            4'd2:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[2][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[2][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[2][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[2][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[2][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[2][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[2][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[2][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[2][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[2][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[2][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[2][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[2][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[2][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[2][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[2][15] ;
                                end
                            4'd3:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[3][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[3][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[3][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[3][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[3][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[3][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[3][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[3][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[3][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[3][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[3][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[3][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[3][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[3][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[3][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[3][15] ;
                                end
                            4'd4:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[4][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[4][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[4][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[4][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[4][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[4][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[4][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[4][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[4][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[4][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[4][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[4][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[4][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[4][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[4][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[4][15] ;
                                end
                            4'd5:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[5][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[5][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[5][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[5][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[5][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[5][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[5][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[5][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[5][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[5][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[5][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[5][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[5][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[5][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[5][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[5][15] ;
                                end
                            4'd6:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[6][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[6][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[6][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[6][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[6][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[6][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[6][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[6][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[6][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[6][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[6][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[6][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[6][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[6][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[6][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[6][15] ;
                                end
                            4'd7:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[7][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[7][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[7][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[7][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[7][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[7][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[7][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[7][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[7][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[7][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[7][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[7][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[7][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[7][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[7][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[7][15] ;
                                end
                            4'd8:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[8][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[8][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[8][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[8][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[8][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[8][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[8][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[8][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[8][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[8][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[8][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[8][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[8][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[8][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[8][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[8][15] ;
                                end
                            4'd9:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[9][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[9][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[9][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[9][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[9][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[9][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[9][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[9][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[9][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[9][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[9][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[9][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[9][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[9][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[9][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[9][15] ;
                                end
                            4'd10:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[10][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[10][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[10][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[10][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[10][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[10][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[10][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[10][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[10][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[10][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[10][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[10][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[10][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[10][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[10][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[10][15] ;
                                end
                            4'd11:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[11][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[11][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[11][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[11][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[11][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[11][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[11][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[11][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[11][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[11][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[11][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[11][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[11][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[11][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[11][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[11][15] ;
                                end
                            4'd12:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[12][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[12][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[12][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[12][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[12][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[12][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[12][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[12][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[12][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[12][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[12][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[12][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[12][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[12][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[12][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[12][15] ;
                                end
                            4'd13:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[13][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[13][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[13][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[13][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[13][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[13][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[13][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[13][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[13][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[13][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[13][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[13][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[13][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[13][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[13][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[13][15] ;
                                end
                            4'd14:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[14][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[14][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[14][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[14][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[14][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[14][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[14][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[14][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[14][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[14][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[14][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[14][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[14][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[14][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[14][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[14][15] ;
                                end
                            4'd15:
                                begin
                                    ROM0_b0     <=  ROM0_st2_arr[15][0]  ;
                                    ROM0_b1     <=  ROM0_st2_arr[15][1]  ;
                                    ROM0_b2     <=  ROM0_st2_arr[15][2]  ;
                                    ROM0_b3     <=  ROM0_st2_arr[15][3]  ;
                                    ROM0_b4     <=  ROM0_st2_arr[15][4]  ;
                                    ROM0_b5     <=  ROM0_st2_arr[15][5]  ;
                                    ROM0_b6     <=  ROM0_st2_arr[15][6]  ;
                                    ROM0_b7     <=  ROM0_st2_arr[15][7]  ;
                                    ROM0_b8     <=  ROM0_st2_arr[15][8]  ;
                                    ROM0_b9     <=  ROM0_st2_arr[15][9]  ;
                                    ROM0_b10    <=  ROM0_st2_arr[15][10] ;
                                    ROM0_b11    <=  ROM0_st2_arr[15][11] ;
                                    ROM0_b12    <=  ROM0_st2_arr[15][12] ;
                                    ROM0_b13    <=  ROM0_st2_arr[15][13] ;
                                    ROM0_b14    <=  ROM0_st2_arr[15][14] ;
                                    ROM0_b15    <=  ROM0_st2_arr[15][15] ;
                                end
                        endcase
                    end
                    2'd3: begin
                        case (MA0)
                            4'd0:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd1:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd2:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd3:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd4:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd5:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd6:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd7:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd8:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd9:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd10:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd11:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd12:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd13:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd14:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                            4'd15:
                                begin
                                    ROM0_b0     <=  ROM0_st3_arr[0]  ;
                                    ROM0_b1     <=  ROM0_st3_arr[1]  ;
                                    ROM0_b2     <=  ROM0_st3_arr[2]  ;
                                    ROM0_b3     <=  ROM0_st3_arr[3]  ;
                                    ROM0_b4     <=  ROM0_st3_arr[4]  ;
                                    ROM0_b5     <=  ROM0_st3_arr[5]  ;
                                    ROM0_b6     <=  ROM0_st3_arr[6]  ;
                                    ROM0_b7     <=  ROM0_st3_arr[7]  ;
                                    ROM0_b8     <=  ROM0_st3_arr[8]  ;
                                    ROM0_b9     <=  ROM0_st3_arr[9]  ;
                                    ROM0_b10    <=  ROM0_st3_arr[10] ;
                                    ROM0_b11    <=  ROM0_st3_arr[11] ;
                                    ROM0_b12    <=  ROM0_st3_arr[12] ;
                                    ROM0_b13    <=  ROM0_st3_arr[13] ;
                                    ROM0_b14    <=  ROM0_st3_arr[14] ;
                                    ROM0_b15    <=  ROM0_st3_arr[15] ;
                                end
                        endcase
                    end
                endcase
            end
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM1_b0     <= 64'd0    ;
            ROM1_b1     <= 64'd0    ;
            ROM1_b2     <= 64'd0    ;
            ROM1_b3     <= 64'd0    ;
            ROM1_b4     <= 64'd0    ;
            ROM1_b5     <= 64'd0    ;
            ROM1_b6     <= 64'd0    ;
            ROM1_b7     <= 64'd0    ;
            ROM1_b8     <= 64'd0    ;
            ROM1_b9     <= 64'd0    ;
            ROM1_b10    <= 64'd0    ;
            ROM1_b11    <= 64'd0    ;
            ROM1_b12    <= 64'd0    ; 
            ROM1_b13    <= 64'd0    ;
            ROM1_b14    <= 64'd0    ; 
            ROM1_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (MA1)
                    4'd0:
                        begin
                            ROM1_b0     <=  ROM1_arr[0][0]  ;
                            ROM1_b1     <=  ROM1_arr[0][1]  ;
                            ROM1_b2     <=  ROM1_arr[0][2]  ;
                            ROM1_b3     <=  ROM1_arr[0][3]  ;
                            ROM1_b4     <=  ROM1_arr[0][4]  ;
                            ROM1_b5     <=  ROM1_arr[0][5]  ;
                            ROM1_b6     <=  ROM1_arr[0][6]  ;
                            ROM1_b7     <=  ROM1_arr[0][7]  ;
                            ROM1_b8     <=  ROM1_arr[0][8]  ;
                            ROM1_b9     <=  ROM1_arr[0][9]  ;
                            ROM1_b10    <=  ROM1_arr[0][10] ;
                            ROM1_b11    <=  ROM1_arr[0][11] ;
                            ROM1_b12    <=  ROM1_arr[0][12] ;
                            ROM1_b13    <=  ROM1_arr[0][13] ;
                            ROM1_b14    <=  ROM1_arr[0][14] ;
                            ROM1_b15    <=  ROM1_arr[0][15] ;
                        end
                    4'd1:
                        begin
                            ROM1_b0     <=  ROM1_arr[1][0]  ;
                            ROM1_b1     <=  ROM1_arr[1][1]  ;
                            ROM1_b2     <=  ROM1_arr[1][2]  ;
                            ROM1_b3     <=  ROM1_arr[1][3]  ;
                            ROM1_b4     <=  ROM1_arr[1][4]  ;
                            ROM1_b5     <=  ROM1_arr[1][5]  ;
                            ROM1_b6     <=  ROM1_arr[1][6]  ;
                            ROM1_b7     <=  ROM1_arr[1][7]  ;
                            ROM1_b8     <=  ROM1_arr[1][8]  ;
                            ROM1_b9     <=  ROM1_arr[1][9]  ;
                            ROM1_b10    <=  ROM1_arr[1][10] ;
                            ROM1_b11    <=  ROM1_arr[1][11] ;
                            ROM1_b12    <=  ROM1_arr[1][12] ;
                            ROM1_b13    <=  ROM1_arr[1][13] ;
                            ROM1_b14    <=  ROM1_arr[1][14] ;
                            ROM1_b15    <=  ROM1_arr[1][15] ;
                        end
                    4'd2:
                        begin
                            ROM1_b0     <=  ROM1_arr[2][0]  ;
                            ROM1_b1     <=  ROM1_arr[2][1]  ;
                            ROM1_b2     <=  ROM1_arr[2][2]  ;
                            ROM1_b3     <=  ROM1_arr[2][3]  ;
                            ROM1_b4     <=  ROM1_arr[2][4]  ;
                            ROM1_b5     <=  ROM1_arr[2][5]  ;
                            ROM1_b6     <=  ROM1_arr[2][6]  ;
                            ROM1_b7     <=  ROM1_arr[2][7]  ;
                            ROM1_b8     <=  ROM1_arr[2][8]  ;
                            ROM1_b9     <=  ROM1_arr[2][9]  ;
                            ROM1_b10    <=  ROM1_arr[2][10] ;
                            ROM1_b11    <=  ROM1_arr[2][11] ;
                            ROM1_b12    <=  ROM1_arr[2][12] ;
                            ROM1_b13    <=  ROM1_arr[2][13] ;
                            ROM1_b14    <=  ROM1_arr[2][14] ;
                            ROM1_b15    <=  ROM1_arr[2][15] ;
                        end
                    4'd3:
                        begin
                            ROM1_b0     <=  ROM1_arr[3][0]  ;
                            ROM1_b1     <=  ROM1_arr[3][1]  ;
                            ROM1_b2     <=  ROM1_arr[3][2]  ;
                            ROM1_b3     <=  ROM1_arr[3][3]  ;
                            ROM1_b4     <=  ROM1_arr[3][4]  ;
                            ROM1_b5     <=  ROM1_arr[3][5]  ;
                            ROM1_b6     <=  ROM1_arr[3][6]  ;
                            ROM1_b7     <=  ROM1_arr[3][7]  ;
                            ROM1_b8     <=  ROM1_arr[3][8]  ;
                            ROM1_b9     <=  ROM1_arr[3][9]  ;
                            ROM1_b10    <=  ROM1_arr[3][10] ;
                            ROM1_b11    <=  ROM1_arr[3][11] ;
                            ROM1_b12    <=  ROM1_arr[3][12] ;
                            ROM1_b13    <=  ROM1_arr[3][13] ;
                            ROM1_b14    <=  ROM1_arr[3][14] ;
                            ROM1_b15    <=  ROM1_arr[3][15] ;
                        end
                    4'd4:
                        begin
                            ROM1_b0     <=  ROM1_arr[4][0]  ;
                            ROM1_b1     <=  ROM1_arr[4][1]  ;
                            ROM1_b2     <=  ROM1_arr[4][2]  ;
                            ROM1_b3     <=  ROM1_arr[4][3]  ;
                            ROM1_b4     <=  ROM1_arr[4][4]  ;
                            ROM1_b5     <=  ROM1_arr[4][5]  ;
                            ROM1_b6     <=  ROM1_arr[4][6]  ;
                            ROM1_b7     <=  ROM1_arr[4][7]  ;
                            ROM1_b8     <=  ROM1_arr[4][8]  ;
                            ROM1_b9     <=  ROM1_arr[4][9]  ;
                            ROM1_b10    <=  ROM1_arr[4][10] ;
                            ROM1_b11    <=  ROM1_arr[4][11] ;
                            ROM1_b12    <=  ROM1_arr[4][12] ;
                            ROM1_b13    <=  ROM1_arr[4][13] ;
                            ROM1_b14    <=  ROM1_arr[4][14] ;
                            ROM1_b15    <=  ROM1_arr[4][15] ;
                        end
                    4'd5:
                        begin
                            ROM1_b0     <=  ROM1_arr[5][0]  ;
                            ROM1_b1     <=  ROM1_arr[5][1]  ;
                            ROM1_b2     <=  ROM1_arr[5][2]  ;
                            ROM1_b3     <=  ROM1_arr[5][3]  ;
                            ROM1_b4     <=  ROM1_arr[5][4]  ;
                            ROM1_b5     <=  ROM1_arr[5][5]  ;
                            ROM1_b6     <=  ROM1_arr[5][6]  ;
                            ROM1_b7     <=  ROM1_arr[5][7]  ;
                            ROM1_b8     <=  ROM1_arr[5][8]  ;
                            ROM1_b9     <=  ROM1_arr[5][9]  ;
                            ROM1_b10    <=  ROM1_arr[5][10] ;
                            ROM1_b11    <=  ROM1_arr[5][11] ;
                            ROM1_b12    <=  ROM1_arr[5][12] ;
                            ROM1_b13    <=  ROM1_arr[5][13] ;
                            ROM1_b14    <=  ROM1_arr[5][14] ;
                            ROM1_b15    <=  ROM1_arr[5][15] ;
                        end
                    4'd6:
                        begin
                            ROM1_b0     <=  ROM1_arr[6][0]  ;
                            ROM1_b1     <=  ROM1_arr[6][1]  ;
                            ROM1_b2     <=  ROM1_arr[6][2]  ;
                            ROM1_b3     <=  ROM1_arr[6][3]  ;
                            ROM1_b4     <=  ROM1_arr[6][4]  ;
                            ROM1_b5     <=  ROM1_arr[6][5]  ;
                            ROM1_b6     <=  ROM1_arr[6][6]  ;
                            ROM1_b7     <=  ROM1_arr[6][7]  ;
                            ROM1_b8     <=  ROM1_arr[6][8]  ;
                            ROM1_b9     <=  ROM1_arr[6][9]  ;
                            ROM1_b10    <=  ROM1_arr[6][10] ;
                            ROM1_b11    <=  ROM1_arr[6][11] ;
                            ROM1_b12    <=  ROM1_arr[6][12] ;
                            ROM1_b13    <=  ROM1_arr[6][13] ;
                            ROM1_b14    <=  ROM1_arr[6][14] ;
                            ROM1_b15    <=  ROM1_arr[6][15] ;
                        end
                    4'd7:
                        begin
                            ROM1_b0     <=  ROM1_arr[7][0]  ;
                            ROM1_b1     <=  ROM1_arr[7][1]  ;
                            ROM1_b2     <=  ROM1_arr[7][2]  ;
                            ROM1_b3     <=  ROM1_arr[7][3]  ;
                            ROM1_b4     <=  ROM1_arr[7][4]  ;
                            ROM1_b5     <=  ROM1_arr[7][5]  ;
                            ROM1_b6     <=  ROM1_arr[7][6]  ;
                            ROM1_b7     <=  ROM1_arr[7][7]  ;
                            ROM1_b8     <=  ROM1_arr[7][8]  ;
                            ROM1_b9     <=  ROM1_arr[7][9]  ;
                            ROM1_b10    <=  ROM1_arr[7][10] ;
                            ROM1_b11    <=  ROM1_arr[7][11] ;
                            ROM1_b12    <=  ROM1_arr[7][12] ;
                            ROM1_b13    <=  ROM1_arr[7][13] ;
                            ROM1_b14    <=  ROM1_arr[7][14] ;
                            ROM1_b15    <=  ROM1_arr[7][15] ;
                        end
                    4'd8:
                        begin
                            ROM1_b0     <=  ROM1_arr[8][0]  ;
                            ROM1_b1     <=  ROM1_arr[8][1]  ;
                            ROM1_b2     <=  ROM1_arr[8][2]  ;
                            ROM1_b3     <=  ROM1_arr[8][3]  ;
                            ROM1_b4     <=  ROM1_arr[8][4]  ;
                            ROM1_b5     <=  ROM1_arr[8][5]  ;
                            ROM1_b6     <=  ROM1_arr[8][6]  ;
                            ROM1_b7     <=  ROM1_arr[8][7]  ;
                            ROM1_b8     <=  ROM1_arr[8][8]  ;
                            ROM1_b9     <=  ROM1_arr[8][9]  ;
                            ROM1_b10    <=  ROM1_arr[8][10] ;
                            ROM1_b11    <=  ROM1_arr[8][11] ;
                            ROM1_b12    <=  ROM1_arr[8][12] ;
                            ROM1_b13    <=  ROM1_arr[8][13] ;
                            ROM1_b14    <=  ROM1_arr[8][14] ;
                            ROM1_b15    <=  ROM1_arr[8][15] ;
                        end
                    4'd9:
                        begin
                            ROM1_b0     <=  ROM1_arr[9][0]  ;
                            ROM1_b1     <=  ROM1_arr[9][1]  ;
                            ROM1_b2     <=  ROM1_arr[9][2]  ;
                            ROM1_b3     <=  ROM1_arr[9][3]  ;
                            ROM1_b4     <=  ROM1_arr[9][4]  ;
                            ROM1_b5     <=  ROM1_arr[9][5]  ;
                            ROM1_b6     <=  ROM1_arr[9][6]  ;
                            ROM1_b7     <=  ROM1_arr[9][7]  ;
                            ROM1_b8     <=  ROM1_arr[9][8]  ;
                            ROM1_b9     <=  ROM1_arr[9][9]  ;
                            ROM1_b10    <=  ROM1_arr[9][10] ;
                            ROM1_b11    <=  ROM1_arr[9][11] ;
                            ROM1_b12    <=  ROM1_arr[9][12] ;
                            ROM1_b13    <=  ROM1_arr[9][13] ;
                            ROM1_b14    <=  ROM1_arr[9][14] ;
                            ROM1_b15    <=  ROM1_arr[9][15] ;
                        end
                    4'd10:
                        begin
                            ROM1_b0     <=  ROM1_arr[10][0]  ;
                            ROM1_b1     <=  ROM1_arr[10][1]  ;
                            ROM1_b2     <=  ROM1_arr[10][2]  ;
                            ROM1_b3     <=  ROM1_arr[10][3]  ;
                            ROM1_b4     <=  ROM1_arr[10][4]  ;
                            ROM1_b5     <=  ROM1_arr[10][5]  ;
                            ROM1_b6     <=  ROM1_arr[10][6]  ;
                            ROM1_b7     <=  ROM1_arr[10][7]  ;
                            ROM1_b8     <=  ROM1_arr[10][8]  ;
                            ROM1_b9     <=  ROM1_arr[10][9]  ;
                            ROM1_b10    <=  ROM1_arr[10][10] ;
                            ROM1_b11    <=  ROM1_arr[10][11] ;
                            ROM1_b12    <=  ROM1_arr[10][12] ;
                            ROM1_b13    <=  ROM1_arr[10][13] ;
                            ROM1_b14    <=  ROM1_arr[10][14] ;
                            ROM1_b15    <=  ROM1_arr[10][15] ;
                        end
                    4'd11:
                        begin
                            ROM1_b0     <=  ROM1_arr[11][0]  ;
                            ROM1_b1     <=  ROM1_arr[11][1]  ;
                            ROM1_b2     <=  ROM1_arr[11][2]  ;
                            ROM1_b3     <=  ROM1_arr[11][3]  ;
                            ROM1_b4     <=  ROM1_arr[11][4]  ;
                            ROM1_b5     <=  ROM1_arr[11][5]  ;
                            ROM1_b6     <=  ROM1_arr[11][6]  ;
                            ROM1_b7     <=  ROM1_arr[11][7]  ;
                            ROM1_b8     <=  ROM1_arr[11][8]  ;
                            ROM1_b9     <=  ROM1_arr[11][9]  ;
                            ROM1_b10    <=  ROM1_arr[11][10] ;
                            ROM1_b11    <=  ROM1_arr[11][11] ;
                            ROM1_b12    <=  ROM1_arr[11][12] ;
                            ROM1_b13    <=  ROM1_arr[11][13] ;
                            ROM1_b14    <=  ROM1_arr[11][14] ;
                            ROM1_b15    <=  ROM1_arr[11][15] ;
                        end
                    4'd12:
                        begin
                            ROM1_b0     <=  ROM1_arr[12][0]  ;
                            ROM1_b1     <=  ROM1_arr[12][1]  ;
                            ROM1_b2     <=  ROM1_arr[12][2]  ;
                            ROM1_b3     <=  ROM1_arr[12][3]  ;
                            ROM1_b4     <=  ROM1_arr[12][4]  ;
                            ROM1_b5     <=  ROM1_arr[12][5]  ;
                            ROM1_b6     <=  ROM1_arr[12][6]  ;
                            ROM1_b7     <=  ROM1_arr[12][7]  ;
                            ROM1_b8     <=  ROM1_arr[12][8]  ;
                            ROM1_b9     <=  ROM1_arr[12][9]  ;
                            ROM1_b10    <=  ROM1_arr[12][10] ;
                            ROM1_b11    <=  ROM1_arr[12][11] ;
                            ROM1_b12    <=  ROM1_arr[12][12] ;
                            ROM1_b13    <=  ROM1_arr[12][13] ;
                            ROM1_b14    <=  ROM1_arr[12][14] ;
                            ROM1_b15    <=  ROM1_arr[12][15] ;
                        end
                    4'd13:
                        begin
                            ROM1_b0     <=  ROM1_arr[13][0]  ;
                            ROM1_b1     <=  ROM1_arr[13][1]  ;
                            ROM1_b2     <=  ROM1_arr[13][2]  ;
                            ROM1_b3     <=  ROM1_arr[13][3]  ;
                            ROM1_b4     <=  ROM1_arr[13][4]  ;
                            ROM1_b5     <=  ROM1_arr[13][5]  ;
                            ROM1_b6     <=  ROM1_arr[13][6]  ;
                            ROM1_b7     <=  ROM1_arr[13][7]  ;
                            ROM1_b8     <=  ROM1_arr[13][8]  ;
                            ROM1_b9     <=  ROM1_arr[13][9]  ;
                            ROM1_b10    <=  ROM1_arr[13][10] ;
                            ROM1_b11    <=  ROM1_arr[13][11] ;
                            ROM1_b12    <=  ROM1_arr[13][12] ;
                            ROM1_b13    <=  ROM1_arr[13][13] ;
                            ROM1_b14    <=  ROM1_arr[13][14] ;
                            ROM1_b15    <=  ROM1_arr[13][15] ;
                        end
                    4'd14:
                        begin
                            ROM1_b0     <=  ROM1_arr[14][0]  ;
                            ROM1_b1     <=  ROM1_arr[14][1]  ;
                            ROM1_b2     <=  ROM1_arr[14][2]  ;
                            ROM1_b3     <=  ROM1_arr[14][3]  ;
                            ROM1_b4     <=  ROM1_arr[14][4]  ;
                            ROM1_b5     <=  ROM1_arr[14][5]  ;
                            ROM1_b6     <=  ROM1_arr[14][6]  ;
                            ROM1_b7     <=  ROM1_arr[14][7]  ;
                            ROM1_b8     <=  ROM1_arr[14][8]  ;
                            ROM1_b9     <=  ROM1_arr[14][9]  ;
                            ROM1_b10    <=  ROM1_arr[14][10] ;
                            ROM1_b11    <=  ROM1_arr[14][11] ;
                            ROM1_b12    <=  ROM1_arr[14][12] ;
                            ROM1_b13    <=  ROM1_arr[14][13] ;
                            ROM1_b14    <=  ROM1_arr[14][14] ;
                            ROM1_b15    <=  ROM1_arr[14][15] ;
                        end
                    4'd15:
                        begin
                            ROM1_b0     <=  ROM1_arr[15][0]  ;
                            ROM1_b1     <=  ROM1_arr[15][1]  ;
                            ROM1_b2     <=  ROM1_arr[15][2]  ;
                            ROM1_b3     <=  ROM1_arr[15][3]  ;
                            ROM1_b4     <=  ROM1_arr[15][4]  ;
                            ROM1_b5     <=  ROM1_arr[15][5]  ;
                            ROM1_b6     <=  ROM1_arr[15][6]  ;
                            ROM1_b7     <=  ROM1_arr[15][7]  ;
                            ROM1_b8     <=  ROM1_arr[15][8]  ;
                            ROM1_b9     <=  ROM1_arr[15][9]  ;
                            ROM1_b10    <=  ROM1_arr[15][10] ;
                            ROM1_b11    <=  ROM1_arr[15][11] ;
                            ROM1_b12    <=  ROM1_arr[15][12] ;
                            ROM1_b13    <=  ROM1_arr[15][13] ;
                            ROM1_b14    <=  ROM1_arr[15][14] ;
                            ROM1_b15    <=  ROM1_arr[15][15] ;
                        end
                endcase
            end
        end
    end

    always @( posedge clk or negedge rst_n ) begin
        if (~rst_n) begin
            ROM2_b0     <= 64'd0    ;
            ROM2_b1     <= 64'd0    ;
            ROM2_b2     <= 64'd0    ;
            ROM2_b3     <= 64'd0    ;
            ROM2_b4     <= 64'd0    ;
            ROM2_b5     <= 64'd0    ;
            ROM2_b6     <= 64'd0    ;
            ROM2_b7     <= 64'd0    ;
            ROM2_b8     <= 64'd0    ;
            ROM2_b9     <= 64'd0    ;
            ROM2_b10    <= 64'd0    ;
            ROM2_b11    <= 64'd0    ;
            ROM2_b12    <= 64'd0    ; 
            ROM2_b13    <= 64'd0    ;
            ROM2_b14    <= 64'd0    ; 
            ROM2_b15    <= 64'd0    ;
        end else begin
            if (~ROM_CEN) begin
                case (MA2)
                    4'd0:
                        begin
                            ROM2_b0     <=  ROM2_arr[0][0]  ;
                            ROM2_b1     <=  ROM2_arr[0][1]  ;
                            ROM2_b2     <=  ROM2_arr[0][2]  ;
                            ROM2_b3     <=  ROM2_arr[0][3]  ;
                            ROM2_b4     <=  ROM2_arr[0][4]  ;
                            ROM2_b5     <=  ROM2_arr[0][5]  ;
                            ROM2_b6     <=  ROM2_arr[0][6]  ;
                            ROM2_b7     <=  ROM2_arr[0][7]  ;
                            ROM2_b8     <=  ROM2_arr[0][8]  ;
                            ROM2_b9     <=  ROM2_arr[0][9]  ;
                            ROM2_b10    <=  ROM2_arr[0][10] ;
                            ROM2_b11    <=  ROM2_arr[0][11] ;
                            ROM2_b12    <=  ROM2_arr[0][12] ;
                            ROM2_b13    <=  ROM2_arr[0][13] ;
                            ROM2_b14    <=  ROM2_arr[0][14] ;
                            ROM2_b15    <=  ROM2_arr[0][15] ;
                        end
                    4'd1:
                        begin
                            ROM2_b0     <=  ROM2_arr[1][0]  ;
                            ROM2_b1     <=  ROM2_arr[1][1]  ;
                            ROM2_b2     <=  ROM2_arr[1][2]  ;
                            ROM2_b3     <=  ROM2_arr[1][3]  ;
                            ROM2_b4     <=  ROM2_arr[1][4]  ;
                            ROM2_b5     <=  ROM2_arr[1][5]  ;
                            ROM2_b6     <=  ROM2_arr[1][6]  ;
                            ROM2_b7     <=  ROM2_arr[1][7]  ;
                            ROM2_b8     <=  ROM2_arr[1][8]  ;
                            ROM2_b9     <=  ROM2_arr[1][9]  ;
                            ROM2_b10    <=  ROM2_arr[1][10] ;
                            ROM2_b11    <=  ROM2_arr[1][11] ;
                            ROM2_b12    <=  ROM2_arr[1][12] ;
                            ROM2_b13    <=  ROM2_arr[1][13] ;
                            ROM2_b14    <=  ROM2_arr[1][14] ;
                            ROM2_b15    <=  ROM2_arr[1][15] ;
                        end
                    4'd2:
                        begin
                            ROM2_b0     <=  ROM2_arr[2][0]  ;
                            ROM2_b1     <=  ROM2_arr[2][1]  ;
                            ROM2_b2     <=  ROM2_arr[2][2]  ;
                            ROM2_b3     <=  ROM2_arr[2][3]  ;
                            ROM2_b4     <=  ROM2_arr[2][4]  ;
                            ROM2_b5     <=  ROM2_arr[2][5]  ;
                            ROM2_b6     <=  ROM2_arr[2][6]  ;
                            ROM2_b7     <=  ROM2_arr[2][7]  ;
                            ROM2_b8     <=  ROM2_arr[2][8]  ;
                            ROM2_b9     <=  ROM2_arr[2][9]  ;
                            ROM2_b10    <=  ROM2_arr[2][10] ;
                            ROM2_b11    <=  ROM2_arr[2][11] ;
                            ROM2_b12    <=  ROM2_arr[2][12] ;
                            ROM2_b13    <=  ROM2_arr[2][13] ;
                            ROM2_b14    <=  ROM2_arr[2][14] ;
                            ROM2_b15    <=  ROM2_arr[2][15] ;
                        end
                    4'd3:
                        begin
                            ROM2_b0     <=  ROM2_arr[3][0]  ;
                            ROM2_b1     <=  ROM2_arr[3][1]  ;
                            ROM2_b2     <=  ROM2_arr[3][2]  ;
                            ROM2_b3     <=  ROM2_arr[3][3]  ;
                            ROM2_b4     <=  ROM2_arr[3][4]  ;
                            ROM2_b5     <=  ROM2_arr[3][5]  ;
                            ROM2_b6     <=  ROM2_arr[3][6]  ;
                            ROM2_b7     <=  ROM2_arr[3][7]  ;
                            ROM2_b8     <=  ROM2_arr[3][8]  ;
                            ROM2_b9     <=  ROM2_arr[3][9]  ;
                            ROM2_b10    <=  ROM2_arr[3][10] ;
                            ROM2_b11    <=  ROM2_arr[3][11] ;
                            ROM2_b12    <=  ROM2_arr[3][12] ;
                            ROM2_b13    <=  ROM2_arr[3][13] ;
                            ROM2_b14    <=  ROM2_arr[3][14] ;
                            ROM2_b15    <=  ROM2_arr[3][15] ;
                        end
                    4'd4:
                        begin
                            ROM2_b0     <=  ROM2_arr[4][0]  ;
                            ROM2_b1     <=  ROM2_arr[4][1]  ;
                            ROM2_b2     <=  ROM2_arr[4][2]  ;
                            ROM2_b3     <=  ROM2_arr[4][3]  ;
                            ROM2_b4     <=  ROM2_arr[4][4]  ;
                            ROM2_b5     <=  ROM2_arr[4][5]  ;
                            ROM2_b6     <=  ROM2_arr[4][6]  ;
                            ROM2_b7     <=  ROM2_arr[4][7]  ;
                            ROM2_b8     <=  ROM2_arr[4][8]  ;
                            ROM2_b9     <=  ROM2_arr[4][9]  ;
                            ROM2_b10    <=  ROM2_arr[4][10] ;
                            ROM2_b11    <=  ROM2_arr[4][11] ;
                            ROM2_b12    <=  ROM2_arr[4][12] ;
                            ROM2_b13    <=  ROM2_arr[4][13] ;
                            ROM2_b14    <=  ROM2_arr[4][14] ;
                            ROM2_b15    <=  ROM2_arr[4][15] ;
                        end
                    4'd5:
                        begin
                            ROM2_b0     <=  ROM2_arr[5][0]  ;
                            ROM2_b1     <=  ROM2_arr[5][1]  ;
                            ROM2_b2     <=  ROM2_arr[5][2]  ;
                            ROM2_b3     <=  ROM2_arr[5][3]  ;
                            ROM2_b4     <=  ROM2_arr[5][4]  ;
                            ROM2_b5     <=  ROM2_arr[5][5]  ;
                            ROM2_b6     <=  ROM2_arr[5][6]  ;
                            ROM2_b7     <=  ROM2_arr[5][7]  ;
                            ROM2_b8     <=  ROM2_arr[5][8]  ;
                            ROM2_b9     <=  ROM2_arr[5][9]  ;
                            ROM2_b10    <=  ROM2_arr[5][10] ;
                            ROM2_b11    <=  ROM2_arr[5][11] ;
                            ROM2_b12    <=  ROM2_arr[5][12] ;
                            ROM2_b13    <=  ROM2_arr[5][13] ;
                            ROM2_b14    <=  ROM2_arr[5][14] ;
                            ROM2_b15    <=  ROM2_arr[5][15] ;
                        end
                    4'd6:
                        begin
                            ROM2_b0     <=  ROM2_arr[6][0]  ;
                            ROM2_b1     <=  ROM2_arr[6][1]  ;
                            ROM2_b2     <=  ROM2_arr[6][2]  ;
                            ROM2_b3     <=  ROM2_arr[6][3]  ;
                            ROM2_b4     <=  ROM2_arr[6][4]  ;
                            ROM2_b5     <=  ROM2_arr[6][5]  ;
                            ROM2_b6     <=  ROM2_arr[6][6]  ;
                            ROM2_b7     <=  ROM2_arr[6][7]  ;
                            ROM2_b8     <=  ROM2_arr[6][8]  ;
                            ROM2_b9     <=  ROM2_arr[6][9]  ;
                            ROM2_b10    <=  ROM2_arr[6][10] ;
                            ROM2_b11    <=  ROM2_arr[6][11] ;
                            ROM2_b12    <=  ROM2_arr[6][12] ;
                            ROM2_b13    <=  ROM2_arr[6][13] ;
                            ROM2_b14    <=  ROM2_arr[6][14] ;
                            ROM2_b15    <=  ROM2_arr[6][15] ;
                        end
                    4'd7:
                        begin
                            ROM2_b0     <=  ROM2_arr[7][0]  ;
                            ROM2_b1     <=  ROM2_arr[7][1]  ;
                            ROM2_b2     <=  ROM2_arr[7][2]  ;
                            ROM2_b3     <=  ROM2_arr[7][3]  ;
                            ROM2_b4     <=  ROM2_arr[7][4]  ;
                            ROM2_b5     <=  ROM2_arr[7][5]  ;
                            ROM2_b6     <=  ROM2_arr[7][6]  ;
                            ROM2_b7     <=  ROM2_arr[7][7]  ;
                            ROM2_b8     <=  ROM2_arr[7][8]  ;
                            ROM2_b9     <=  ROM2_arr[7][9]  ;
                            ROM2_b10    <=  ROM2_arr[7][10] ;
                            ROM2_b11    <=  ROM2_arr[7][11] ;
                            ROM2_b12    <=  ROM2_arr[7][12] ;
                            ROM2_b13    <=  ROM2_arr[7][13] ;
                            ROM2_b14    <=  ROM2_arr[7][14] ;
                            ROM2_b15    <=  ROM2_arr[7][15] ;
                        end
                    4'd8:
                        begin
                            ROM2_b0     <=  ROM2_arr[8][0]  ;
                            ROM2_b1     <=  ROM2_arr[8][1]  ;
                            ROM2_b2     <=  ROM2_arr[8][2]  ;
                            ROM2_b3     <=  ROM2_arr[8][3]  ;
                            ROM2_b4     <=  ROM2_arr[8][4]  ;
                            ROM2_b5     <=  ROM2_arr[8][5]  ;
                            ROM2_b6     <=  ROM2_arr[8][6]  ;
                            ROM2_b7     <=  ROM2_arr[8][7]  ;
                            ROM2_b8     <=  ROM2_arr[8][8]  ;
                            ROM2_b9     <=  ROM2_arr[8][9]  ;
                            ROM2_b10    <=  ROM2_arr[8][10] ;
                            ROM2_b11    <=  ROM2_arr[8][11] ;
                            ROM2_b12    <=  ROM2_arr[8][12] ;
                            ROM2_b13    <=  ROM2_arr[8][13] ;
                            ROM2_b14    <=  ROM2_arr[8][14] ;
                            ROM2_b15    <=  ROM2_arr[8][15] ;
                        end
                    4'd9:
                        begin
                            ROM2_b0     <=  ROM2_arr[9][0]  ;
                            ROM2_b1     <=  ROM2_arr[9][1]  ;
                            ROM2_b2     <=  ROM2_arr[9][2]  ;
                            ROM2_b3     <=  ROM2_arr[9][3]  ;
                            ROM2_b4     <=  ROM2_arr[9][4]  ;
                            ROM2_b5     <=  ROM2_arr[9][5]  ;
                            ROM2_b6     <=  ROM2_arr[9][6]  ;
                            ROM2_b7     <=  ROM2_arr[9][7]  ;
                            ROM2_b8     <=  ROM2_arr[9][8]  ;
                            ROM2_b9     <=  ROM2_arr[9][9]  ;
                            ROM2_b10    <=  ROM2_arr[9][10] ;
                            ROM2_b11    <=  ROM2_arr[9][11] ;
                            ROM2_b12    <=  ROM2_arr[9][12] ;
                            ROM2_b13    <=  ROM2_arr[9][13] ;
                            ROM2_b14    <=  ROM2_arr[9][14] ;
                            ROM2_b15    <=  ROM2_arr[9][15] ;
                        end
                    4'd10:
                        begin
                            ROM2_b0     <=  ROM2_arr[10][0]  ;
                            ROM2_b1     <=  ROM2_arr[10][1]  ;
                            ROM2_b2     <=  ROM2_arr[10][2]  ;
                            ROM2_b3     <=  ROM2_arr[10][3]  ;
                            ROM2_b4     <=  ROM2_arr[10][4]  ;
                            ROM2_b5     <=  ROM2_arr[10][5]  ;
                            ROM2_b6     <=  ROM2_arr[10][6]  ;
                            ROM2_b7     <=  ROM2_arr[10][7]  ;
                            ROM2_b8     <=  ROM2_arr[10][8]  ;
                            ROM2_b9     <=  ROM2_arr[10][9]  ;
                            ROM2_b10    <=  ROM2_arr[10][10] ;
                            ROM2_b11    <=  ROM2_arr[10][11] ;
                            ROM2_b12    <=  ROM2_arr[10][12] ;
                            ROM2_b13    <=  ROM2_arr[10][13] ;
                            ROM2_b14    <=  ROM2_arr[10][14] ;
                            ROM2_b15    <=  ROM2_arr[10][15] ;
                        end
                    4'd11:
                        begin
                            ROM2_b0     <=  ROM2_arr[11][0]  ;
                            ROM2_b1     <=  ROM2_arr[11][1]  ;
                            ROM2_b2     <=  ROM2_arr[11][2]  ;
                            ROM2_b3     <=  ROM2_arr[11][3]  ;
                            ROM2_b4     <=  ROM2_arr[11][4]  ;
                            ROM2_b5     <=  ROM2_arr[11][5]  ;
                            ROM2_b6     <=  ROM2_arr[11][6]  ;
                            ROM2_b7     <=  ROM2_arr[11][7]  ;
                            ROM2_b8     <=  ROM2_arr[11][8]  ;
                            ROM2_b9     <=  ROM2_arr[11][9]  ;
                            ROM2_b10    <=  ROM2_arr[11][10] ;
                            ROM2_b11    <=  ROM2_arr[11][11] ;
                            ROM2_b12    <=  ROM2_arr[11][12] ;
                            ROM2_b13    <=  ROM2_arr[11][13] ;
                            ROM2_b14    <=  ROM2_arr[11][14] ;
                            ROM2_b15    <=  ROM2_arr[11][15] ;
                        end
                    4'd12:
                        begin
                            ROM2_b0     <=  ROM2_arr[12][0]  ;
                            ROM2_b1     <=  ROM2_arr[12][1]  ;
                            ROM2_b2     <=  ROM2_arr[12][2]  ;
                            ROM2_b3     <=  ROM2_arr[12][3]  ;
                            ROM2_b4     <=  ROM2_arr[12][4]  ;
                            ROM2_b5     <=  ROM2_arr[12][5]  ;
                            ROM2_b6     <=  ROM2_arr[12][6]  ;
                            ROM2_b7     <=  ROM2_arr[12][7]  ;
                            ROM2_b8     <=  ROM2_arr[12][8]  ;
                            ROM2_b9     <=  ROM2_arr[12][9]  ;
                            ROM2_b10    <=  ROM2_arr[12][10] ;
                            ROM2_b11    <=  ROM2_arr[12][11] ;
                            ROM2_b12    <=  ROM2_arr[12][12] ;
                            ROM2_b13    <=  ROM2_arr[12][13] ;
                            ROM2_b14    <=  ROM2_arr[12][14] ;
                            ROM2_b15    <=  ROM2_arr[12][15] ;
                        end
                    4'd13:
                        begin
                            ROM2_b0     <=  ROM2_arr[13][0]  ;
                            ROM2_b1     <=  ROM2_arr[13][1]  ;
                            ROM2_b2     <=  ROM2_arr[13][2]  ;
                            ROM2_b3     <=  ROM2_arr[13][3]  ;
                            ROM2_b4     <=  ROM2_arr[13][4]  ;
                            ROM2_b5     <=  ROM2_arr[13][5]  ;
                            ROM2_b6     <=  ROM2_arr[13][6]  ;
                            ROM2_b7     <=  ROM2_arr[13][7]  ;
                            ROM2_b8     <=  ROM2_arr[13][8]  ;
                            ROM2_b9     <=  ROM2_arr[13][9]  ;
                            ROM2_b10    <=  ROM2_arr[13][10] ;
                            ROM2_b11    <=  ROM2_arr[13][11] ;
                            ROM2_b12    <=  ROM2_arr[13][12] ;
                            ROM2_b13    <=  ROM2_arr[13][13] ;
                            ROM2_b14    <=  ROM2_arr[13][14] ;
                            ROM2_b15    <=  ROM2_arr[13][15] ;
                        end
                    4'd14:
                        begin
                            ROM2_b0     <=  ROM2_arr[14][0]  ;
                            ROM2_b1     <=  ROM2_arr[14][1]  ;
                            ROM2_b2     <=  ROM2_arr[14][2]  ;
                            ROM2_b3     <=  ROM2_arr[14][3]  ;
                            ROM2_b4     <=  ROM2_arr[14][4]  ;
                            ROM2_b5     <=  ROM2_arr[14][5]  ;
                            ROM2_b6     <=  ROM2_arr[14][6]  ;
                            ROM2_b7     <=  ROM2_arr[14][7]  ;
                            ROM2_b8     <=  ROM2_arr[14][8]  ;
                            ROM2_b9     <=  ROM2_arr[14][9]  ;
                            ROM2_b10    <=  ROM2_arr[14][10] ;
                            ROM2_b11    <=  ROM2_arr[14][11] ;
                            ROM2_b12    <=  ROM2_arr[14][12] ;
                            ROM2_b13    <=  ROM2_arr[14][13] ;
                            ROM2_b14    <=  ROM2_arr[14][14] ;
                            ROM2_b15    <=  ROM2_arr[14][15] ;
                        end
                    4'd15:
                        begin
                            ROM2_b0     <=  ROM2_arr[15][0]  ;
                            ROM2_b1     <=  ROM2_arr[15][1]  ;
                            ROM2_b2     <=  ROM2_arr[15][2]  ;
                            ROM2_b3     <=  ROM2_arr[15][3]  ;
                            ROM2_b4     <=  ROM2_arr[15][4]  ;
                            ROM2_b5     <=  ROM2_arr[15][5]  ;
                            ROM2_b6     <=  ROM2_arr[15][6]  ;
                            ROM2_b7     <=  ROM2_arr[15][7]  ;
                            ROM2_b8     <=  ROM2_arr[15][8]  ;
                            ROM2_b9     <=  ROM2_arr[15][9]  ;
                            ROM2_b10    <=  ROM2_arr[15][10] ;
                            ROM2_b11    <=  ROM2_arr[15][11] ;
                            ROM2_b12    <=  ROM2_arr[15][12] ;
                            ROM2_b13    <=  ROM2_arr[15][13] ;
                            ROM2_b14    <=  ROM2_arr[15][14] ;
                            ROM2_b15    <=  ROM2_arr[15][15] ;
                        end
                endcase
            end
        end
    end
endmodule